-- generated with romgen by MikeJ
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity BBC_BASIC_ROM is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of BBC_BASIC_ROM is


  type ROM_ARRAY is array(0 to 16383) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"C9",x"01",x"F0",x"1F",x"60",x"EA",x"60",x"0E", -- 0x0000
    x"01",x"42",x"41",x"53",x"49",x"43",x"00",x"28", -- 0x0008
    x"43",x"29",x"31",x"39",x"38",x"32",x"20",x"41", -- 0x0010
    x"63",x"6F",x"72",x"6E",x"0A",x"0D",x"00",x"00", -- 0x0018
    x"80",x"00",x"00",x"A9",x"84",x"20",x"F4",x"FF", -- 0x0020
    x"86",x"06",x"84",x"07",x"A9",x"83",x"20",x"F4", -- 0x0028
    x"FF",x"84",x"18",x"A2",x"00",x"86",x"1F",x"8E", -- 0x0030
    x"02",x"04",x"8E",x"03",x"04",x"CA",x"86",x"23", -- 0x0038
    x"A2",x"0A",x"8E",x"00",x"04",x"CA",x"8E",x"01", -- 0x0040
    x"04",x"A9",x"01",x"25",x"11",x"05",x"0D",x"05", -- 0x0048
    x"0E",x"05",x"0F",x"05",x"10",x"D0",x"0C",x"A9", -- 0x0050
    x"41",x"85",x"0D",x"A9",x"52",x"85",x"0E",x"A9", -- 0x0058
    x"57",x"85",x"0F",x"A9",x"02",x"8D",x"02",x"02", -- 0x0060
    x"A9",x"B4",x"8D",x"03",x"02",x"58",x"4C",x"DD", -- 0x0068
    x"8A",x"41",x"4E",x"44",x"80",x"00",x"41",x"42", -- 0x0070
    x"53",x"94",x"00",x"41",x"43",x"53",x"95",x"00", -- 0x0078
    x"41",x"44",x"56",x"41",x"4C",x"96",x"00",x"41", -- 0x0080
    x"53",x"43",x"97",x"00",x"41",x"53",x"4E",x"98", -- 0x0088
    x"00",x"41",x"54",x"4E",x"99",x"00",x"41",x"55", -- 0x0090
    x"54",x"4F",x"C6",x"10",x"42",x"47",x"45",x"54", -- 0x0098
    x"9A",x"01",x"42",x"50",x"55",x"54",x"D5",x"03", -- 0x00A0
    x"43",x"4F",x"4C",x"4F",x"55",x"52",x"FB",x"02", -- 0x00A8
    x"43",x"41",x"4C",x"4C",x"D6",x"02",x"43",x"48", -- 0x00B0
    x"41",x"49",x"4E",x"D7",x"02",x"43",x"48",x"52", -- 0x00B8
    x"24",x"BD",x"00",x"43",x"4C",x"45",x"41",x"52", -- 0x00C0
    x"D8",x"01",x"43",x"4C",x"4F",x"53",x"45",x"D9", -- 0x00C8
    x"03",x"43",x"4C",x"47",x"DA",x"01",x"43",x"4C", -- 0x00D0
    x"53",x"DB",x"01",x"43",x"4F",x"53",x"9B",x"00", -- 0x00D8
    x"43",x"4F",x"55",x"4E",x"54",x"9C",x"01",x"44", -- 0x00E0
    x"41",x"54",x"41",x"DC",x"20",x"44",x"45",x"47", -- 0x00E8
    x"9D",x"00",x"44",x"45",x"46",x"DD",x"00",x"44", -- 0x00F0
    x"45",x"4C",x"45",x"54",x"45",x"C7",x"10",x"44", -- 0x00F8
    x"49",x"56",x"81",x"00",x"44",x"49",x"4D",x"DE", -- 0x0100
    x"02",x"44",x"52",x"41",x"57",x"DF",x"02",x"45", -- 0x0108
    x"4E",x"44",x"50",x"52",x"4F",x"43",x"E1",x"01", -- 0x0110
    x"45",x"4E",x"44",x"E0",x"01",x"45",x"4E",x"56", -- 0x0118
    x"45",x"4C",x"4F",x"50",x"45",x"E2",x"02",x"45", -- 0x0120
    x"4C",x"53",x"45",x"8B",x"14",x"45",x"56",x"41", -- 0x0128
    x"4C",x"A0",x"00",x"45",x"52",x"4C",x"9E",x"01", -- 0x0130
    x"45",x"52",x"52",x"4F",x"52",x"85",x"04",x"45", -- 0x0138
    x"4F",x"46",x"C5",x"01",x"45",x"4F",x"52",x"82", -- 0x0140
    x"00",x"45",x"52",x"52",x"9F",x"01",x"45",x"58", -- 0x0148
    x"50",x"A1",x"00",x"45",x"58",x"54",x"A2",x"01", -- 0x0150
    x"46",x"4F",x"52",x"E3",x"02",x"46",x"41",x"4C", -- 0x0158
    x"53",x"45",x"A3",x"01",x"46",x"4E",x"A4",x"08", -- 0x0160
    x"47",x"4F",x"54",x"4F",x"E5",x"12",x"47",x"45", -- 0x0168
    x"54",x"24",x"BE",x"00",x"47",x"45",x"54",x"A5", -- 0x0170
    x"00",x"47",x"4F",x"53",x"55",x"42",x"E4",x"12", -- 0x0178
    x"47",x"43",x"4F",x"4C",x"E6",x"02",x"48",x"49", -- 0x0180
    x"4D",x"45",x"4D",x"93",x"43",x"49",x"4E",x"50", -- 0x0188
    x"55",x"54",x"E8",x"02",x"49",x"46",x"E7",x"02", -- 0x0190
    x"49",x"4E",x"4B",x"45",x"59",x"24",x"BF",x"00", -- 0x0198
    x"49",x"4E",x"4B",x"45",x"59",x"A6",x"00",x"49", -- 0x01A0
    x"4E",x"54",x"A8",x"00",x"49",x"4E",x"53",x"54", -- 0x01A8
    x"52",x"28",x"A7",x"00",x"4C",x"49",x"53",x"54", -- 0x01B0
    x"C9",x"10",x"4C",x"49",x"4E",x"45",x"86",x"00", -- 0x01B8
    x"4C",x"4F",x"41",x"44",x"C8",x"02",x"4C",x"4F", -- 0x01C0
    x"4D",x"45",x"4D",x"92",x"43",x"4C",x"4F",x"43", -- 0x01C8
    x"41",x"4C",x"EA",x"02",x"4C",x"45",x"46",x"54", -- 0x01D0
    x"24",x"28",x"C0",x"00",x"4C",x"45",x"4E",x"A9", -- 0x01D8
    x"00",x"4C",x"45",x"54",x"E9",x"04",x"4C",x"4F", -- 0x01E0
    x"47",x"AB",x"00",x"4C",x"4E",x"AA",x"00",x"4D", -- 0x01E8
    x"49",x"44",x"24",x"28",x"C1",x"00",x"4D",x"4F", -- 0x01F0
    x"44",x"45",x"EB",x"02",x"4D",x"4F",x"44",x"83", -- 0x01F8
    x"00",x"4D",x"4F",x"56",x"45",x"EC",x"02",x"4E", -- 0x0200
    x"45",x"58",x"54",x"ED",x"02",x"4E",x"45",x"57", -- 0x0208
    x"CA",x"01",x"4E",x"4F",x"54",x"AC",x"00",x"4F", -- 0x0210
    x"4C",x"44",x"CB",x"01",x"4F",x"4E",x"EE",x"02", -- 0x0218
    x"4F",x"46",x"46",x"87",x"00",x"4F",x"52",x"84", -- 0x0220
    x"00",x"4F",x"50",x"45",x"4E",x"49",x"4E",x"8E", -- 0x0228
    x"00",x"4F",x"50",x"45",x"4E",x"4F",x"55",x"54", -- 0x0230
    x"AE",x"00",x"4F",x"50",x"45",x"4E",x"55",x"50", -- 0x0238
    x"AD",x"00",x"4F",x"53",x"43",x"4C",x"49",x"FF", -- 0x0240
    x"02",x"50",x"52",x"49",x"4E",x"54",x"F1",x"02", -- 0x0248
    x"50",x"41",x"47",x"45",x"90",x"43",x"50",x"54", -- 0x0250
    x"52",x"8F",x"43",x"50",x"49",x"AF",x"01",x"50", -- 0x0258
    x"4C",x"4F",x"54",x"F0",x"02",x"50",x"4F",x"49", -- 0x0260
    x"4E",x"54",x"28",x"B0",x"00",x"50",x"52",x"4F", -- 0x0268
    x"43",x"F2",x"0A",x"50",x"4F",x"53",x"B1",x"01", -- 0x0270
    x"52",x"45",x"54",x"55",x"52",x"4E",x"F8",x"01", -- 0x0278
    x"52",x"45",x"50",x"45",x"41",x"54",x"F5",x"00", -- 0x0280
    x"52",x"45",x"50",x"4F",x"52",x"54",x"F6",x"01", -- 0x0288
    x"52",x"45",x"41",x"44",x"F3",x"02",x"52",x"45", -- 0x0290
    x"4D",x"F4",x"20",x"52",x"55",x"4E",x"F9",x"01", -- 0x0298
    x"52",x"41",x"44",x"B2",x"00",x"52",x"45",x"53", -- 0x02A0
    x"54",x"4F",x"52",x"45",x"F7",x"12",x"52",x"49", -- 0x02A8
    x"47",x"48",x"54",x"24",x"28",x"C2",x"00",x"52", -- 0x02B0
    x"4E",x"44",x"B3",x"01",x"52",x"45",x"4E",x"55", -- 0x02B8
    x"4D",x"42",x"45",x"52",x"CC",x"10",x"53",x"54", -- 0x02C0
    x"45",x"50",x"88",x"00",x"53",x"41",x"56",x"45", -- 0x02C8
    x"CD",x"02",x"53",x"47",x"4E",x"B4",x"00",x"53", -- 0x02D0
    x"49",x"4E",x"B5",x"00",x"53",x"51",x"52",x"B6", -- 0x02D8
    x"00",x"53",x"50",x"43",x"89",x"00",x"53",x"54", -- 0x02E0
    x"52",x"24",x"C3",x"00",x"53",x"54",x"52",x"49", -- 0x02E8
    x"4E",x"47",x"24",x"28",x"C4",x"00",x"53",x"4F", -- 0x02F0
    x"55",x"4E",x"44",x"D4",x"02",x"53",x"54",x"4F", -- 0x02F8
    x"50",x"FA",x"01",x"54",x"41",x"4E",x"B7",x"00", -- 0x0300
    x"54",x"48",x"45",x"4E",x"8C",x"14",x"54",x"4F", -- 0x0308
    x"B8",x"00",x"54",x"41",x"42",x"28",x"8A",x"00", -- 0x0310
    x"54",x"52",x"41",x"43",x"45",x"FC",x"12",x"54", -- 0x0318
    x"49",x"4D",x"45",x"91",x"43",x"54",x"52",x"55", -- 0x0320
    x"45",x"B9",x"01",x"55",x"4E",x"54",x"49",x"4C", -- 0x0328
    x"FD",x"02",x"55",x"53",x"52",x"BA",x"00",x"56", -- 0x0330
    x"44",x"55",x"EF",x"02",x"56",x"41",x"4C",x"BB", -- 0x0338
    x"00",x"56",x"50",x"4F",x"53",x"BC",x"01",x"57", -- 0x0340
    x"49",x"44",x"54",x"48",x"FE",x"02",x"50",x"41", -- 0x0348
    x"47",x"45",x"D0",x"00",x"50",x"54",x"52",x"CF", -- 0x0350
    x"00",x"54",x"49",x"4D",x"45",x"D1",x"00",x"4C", -- 0x0358
    x"4F",x"4D",x"45",x"4D",x"D2",x"00",x"48",x"49", -- 0x0360
    x"4D",x"45",x"4D",x"D3",x"00",x"78",x"47",x"C0", -- 0x0368
    x"B4",x"FC",x"03",x"6A",x"D4",x"33",x"9E",x"DA", -- 0x0370
    x"07",x"6F",x"8D",x"F7",x"C2",x"9F",x"A6",x"E9", -- 0x0378
    x"91",x"46",x"CA",x"95",x"B9",x"AD",x"E2",x"78", -- 0x0380
    x"D1",x"FE",x"A8",x"D1",x"80",x"7C",x"CB",x"41", -- 0x0388
    x"6D",x"B1",x"49",x"88",x"98",x"B4",x"BE",x"DC", -- 0x0390
    x"C4",x"D2",x"2F",x"76",x"BD",x"BF",x"26",x"CC", -- 0x0398
    x"39",x"EE",x"94",x"C2",x"B8",x"AC",x"31",x"24", -- 0x03A0
    x"9C",x"DA",x"B6",x"A3",x"F3",x"2A",x"30",x"83", -- 0x03A8
    x"C9",x"6F",x"5D",x"4C",x"58",x"D2",x"2A",x"8D", -- 0x03B0
    x"99",x"BD",x"C4",x"7D",x"7D",x"2F",x"E8",x"C8", -- 0x03B8
    x"56",x"72",x"C4",x"88",x"CC",x"7A",x"C2",x"44", -- 0x03C0
    x"E4",x"23",x"9A",x"E4",x"95",x"15",x"2F",x"F1", -- 0x03C8
    x"9A",x"04",x"1F",x"7D",x"E4",x"E4",x"E6",x"B6", -- 0x03D0
    x"11",x"D0",x"8E",x"95",x"B1",x"A0",x"C2",x"BF", -- 0x03D8
    x"BF",x"AE",x"AE",x"AE",x"AF",x"AD",x"A8",x"AB", -- 0x03E0
    x"AC",x"A8",x"A9",x"BF",x"A9",x"AE",x"AB",x"AF", -- 0x03E8
    x"AF",x"AB",x"AA",x"BF",x"AE",x"B1",x"AF",x"AC", -- 0x03F0
    x"AC",x"AC",x"AE",x"A7",x"AB",x"AC",x"BF",x"BF", -- 0x03F8
    x"AB",x"AB",x"AB",x"AB",x"AF",x"AB",x"A9",x"A7", -- 0x0400
    x"A6",x"AE",x"AC",x"AB",x"AC",x"AB",x"B3",x"AF", -- 0x0408
    x"B0",x"AF",x"B0",x"AF",x"B0",x"B0",x"AC",x"90", -- 0x0410
    x"8F",x"BF",x"B5",x"8A",x"8A",x"8F",x"BE",x"98", -- 0x0418
    x"BF",x"92",x"92",x"92",x"92",x"B4",x"BF",x"8E", -- 0x0420
    x"BF",x"92",x"BF",x"8E",x"8E",x"8B",x"8B",x"91", -- 0x0428
    x"93",x"8A",x"93",x"B4",x"B7",x"B8",x"B8",x"93", -- 0x0430
    x"98",x"BA",x"8B",x"93",x"93",x"93",x"B6",x"B9", -- 0x0438
    x"94",x"93",x"8D",x"93",x"BB",x"8B",x"BB",x"BF", -- 0x0440
    x"BA",x"B8",x"BD",x"8A",x"93",x"92",x"BB",x"B4", -- 0x0448
    x"BE",x"4B",x"83",x"84",x"89",x"96",x"B8",x"B9", -- 0x0450
    x"D8",x"D9",x"F0",x"01",x"10",x"81",x"90",x"89", -- 0x0458
    x"93",x"A3",x"A4",x"A9",x"38",x"39",x"78",x"01", -- 0x0460
    x"13",x"21",x"63",x"73",x"B1",x"A9",x"C5",x"0C", -- 0x0468
    x"C3",x"D3",x"C4",x"F2",x"41",x"83",x"B0",x"81", -- 0x0470
    x"43",x"6C",x"72",x"EC",x"F2",x"A3",x"C3",x"18", -- 0x0478
    x"19",x"34",x"B0",x"72",x"98",x"99",x"81",x"98", -- 0x0480
    x"99",x"14",x"35",x"0A",x"0D",x"0D",x"0D",x"0D", -- 0x0488
    x"10",x"10",x"25",x"25",x"39",x"41",x"41",x"41", -- 0x0490
    x"41",x"4A",x"4A",x"4C",x"4C",x"4C",x"50",x"50", -- 0x0498
    x"52",x"53",x"53",x"53",x"08",x"08",x"08",x"09", -- 0x04A0
    x"09",x"0A",x"0A",x"0A",x"05",x"15",x"3E",x"04", -- 0x04A8
    x"0D",x"30",x"4C",x"06",x"32",x"49",x"49",x"10", -- 0x04B0
    x"25",x"0E",x"0E",x"09",x"29",x"2A",x"30",x"30", -- 0x04B8
    x"4E",x"4E",x"4E",x"3E",x"16",x"00",x"18",x"D8", -- 0x04C0
    x"58",x"B8",x"CA",x"88",x"E8",x"C8",x"EA",x"48", -- 0x04C8
    x"08",x"68",x"28",x"40",x"60",x"38",x"F8",x"78", -- 0x04D0
    x"AA",x"A8",x"BA",x"8A",x"9A",x"98",x"90",x"B0", -- 0x04D8
    x"F0",x"30",x"D0",x"10",x"50",x"70",x"21",x"41", -- 0x04E0
    x"01",x"61",x"C1",x"A1",x"E1",x"06",x"46",x"26", -- 0x04E8
    x"66",x"C6",x"E6",x"E0",x"C0",x"20",x"4C",x"20", -- 0x04F0
    x"A2",x"A0",x"81",x"86",x"84",x"A9",x"FF",x"85", -- 0x04F8
    x"28",x"4C",x"A3",x"8B",x"A9",x"03",x"85",x"28", -- 0x0500
    x"20",x"97",x"8A",x"C9",x"5D",x"F0",x"EE",x"20", -- 0x0508
    x"6D",x"98",x"C6",x"0A",x"20",x"BA",x"85",x"C6", -- 0x0510
    x"0A",x"A5",x"28",x"4A",x"90",x"60",x"A5",x"1E", -- 0x0518
    x"69",x"04",x"85",x"3F",x"A5",x"38",x"20",x"45", -- 0x0520
    x"B5",x"A5",x"37",x"20",x"62",x"B5",x"A2",x"FC", -- 0x0528
    x"A4",x"39",x"10",x"02",x"A4",x"36",x"84",x"38", -- 0x0530
    x"F0",x"1C",x"A0",x"00",x"E8",x"D0",x"0D",x"20", -- 0x0538
    x"25",x"BC",x"A6",x"3F",x"20",x"65",x"B5",x"CA", -- 0x0540
    x"D0",x"FA",x"A2",x"FD",x"B1",x"3A",x"20",x"62", -- 0x0548
    x"B5",x"C8",x"C6",x"38",x"D0",x"E6",x"E8",x"10", -- 0x0550
    x"0C",x"20",x"65",x"B5",x"20",x"58",x"B5",x"20", -- 0x0558
    x"58",x"B5",x"4C",x"56",x"85",x"A0",x"00",x"B1", -- 0x0560
    x"0B",x"C9",x"3A",x"F0",x"0A",x"C9",x"0D",x"F0", -- 0x0568
    x"0A",x"20",x"0E",x"B5",x"C8",x"D0",x"F0",x"C4", -- 0x0570
    x"0A",x"90",x"F6",x"20",x"25",x"BC",x"A4",x"0A", -- 0x0578
    x"88",x"C8",x"B1",x"0B",x"C9",x"3A",x"F0",x"04", -- 0x0580
    x"C9",x"0D",x"D0",x"F5",x"20",x"59",x"98",x"88", -- 0x0588
    x"B1",x"0B",x"C9",x"3A",x"F0",x"0C",x"A5",x"0C", -- 0x0590
    x"C9",x"07",x"D0",x"03",x"4C",x"F6",x"8A",x"20", -- 0x0598
    x"90",x"98",x"4C",x"08",x"85",x"20",x"82",x"95", -- 0x05A0
    x"F0",x"5A",x"B0",x"58",x"20",x"94",x"BD",x"20", -- 0x05A8
    x"3A",x"AE",x"85",x"27",x"20",x"B4",x"B4",x"20", -- 0x05B0
    x"27",x"88",x"A2",x"03",x"20",x"97",x"8A",x"A0", -- 0x05B8
    x"00",x"84",x"3D",x"C9",x"3A",x"F0",x"64",x"C9", -- 0x05C0
    x"0D",x"F0",x"60",x"C9",x"5C",x"F0",x"5C",x"C9", -- 0x05C8
    x"2E",x"F0",x"D2",x"C6",x"0A",x"A4",x"0A",x"E6", -- 0x05D0
    x"0A",x"B1",x"0B",x"30",x"2A",x"C9",x"20",x"F0", -- 0x05D8
    x"10",x"A0",x"05",x"0A",x"0A",x"0A",x"0A",x"26", -- 0x05E0
    x"3D",x"26",x"3E",x"88",x"D0",x"F8",x"CA",x"D0", -- 0x05E8
    x"E4",x"A2",x"3A",x"A5",x"3D",x"DD",x"50",x"84", -- 0x05F0
    x"D0",x"07",x"BC",x"8A",x"84",x"C4",x"3E",x"F0", -- 0x05F8
    x"1F",x"CA",x"D0",x"F1",x"4C",x"2A",x"98",x"A2", -- 0x0600
    x"22",x"C9",x"80",x"F0",x"13",x"E8",x"C9",x"82", -- 0x0608
    x"F0",x"0E",x"E8",x"C9",x"84",x"D0",x"ED",x"E6", -- 0x0610
    x"0A",x"C8",x"B1",x"0B",x"C9",x"41",x"D0",x"E4", -- 0x0618
    x"BD",x"C4",x"84",x"85",x"29",x"A0",x"01",x"E0", -- 0x0620
    x"1A",x"B0",x"48",x"AD",x"40",x"04",x"85",x"37", -- 0x0628
    x"84",x"39",x"A6",x"28",x"E0",x"04",x"AE",x"41", -- 0x0630
    x"04",x"86",x"38",x"90",x"06",x"AD",x"3C",x"04", -- 0x0638
    x"AE",x"3D",x"04",x"85",x"3A",x"86",x"3B",x"98", -- 0x0640
    x"F0",x"28",x"10",x"04",x"A4",x"36",x"F0",x"22", -- 0x0648
    x"88",x"B9",x"29",x"00",x"24",x"39",x"10",x"03", -- 0x0650
    x"B9",x"00",x"06",x"91",x"3A",x"EE",x"40",x"04", -- 0x0658
    x"D0",x"03",x"EE",x"41",x"04",x"90",x"08",x"EE", -- 0x0660
    x"3C",x"04",x"D0",x"03",x"EE",x"3D",x"04",x"98", -- 0x0668
    x"D0",x"DE",x"60",x"E0",x"22",x"B0",x"40",x"20", -- 0x0670
    x"21",x"88",x"18",x"A5",x"2A",x"ED",x"40",x"04", -- 0x0678
    x"A8",x"A5",x"2B",x"ED",x"41",x"04",x"C0",x"01", -- 0x0680
    x"88",x"E9",x"00",x"F0",x"25",x"C9",x"FF",x"F0", -- 0x0688
    x"1C",x"A5",x"28",x"4A",x"F0",x"0F",x"00",x"01", -- 0x0690
    x"4F",x"75",x"74",x"20",x"6F",x"66",x"20",x"72", -- 0x0698
    x"61",x"6E",x"67",x"65",x"00",x"A8",x"84",x"2A", -- 0x06A0
    x"A0",x"02",x"4C",x"2B",x"86",x"98",x"30",x"F6", -- 0x06A8
    x"10",x"DF",x"98",x"10",x"F1",x"30",x"DA",x"E0", -- 0x06B0
    x"29",x"B0",x"18",x"20",x"97",x"8A",x"C9",x"23", -- 0x06B8
    x"D0",x"18",x"20",x"2F",x"88",x"20",x"21",x"88", -- 0x06C0
    x"A5",x"2B",x"F0",x"DC",x"00",x"02",x"42",x"79", -- 0x06C8
    x"74",x"65",x"00",x"E0",x"36",x"D0",x"68",x"20", -- 0x06D0
    x"97",x"8A",x"C9",x"28",x"D0",x"37",x"20",x"21", -- 0x06D8
    x"88",x"20",x"97",x"8A",x"C9",x"29",x"D0",x"13", -- 0x06E0
    x"20",x"97",x"8A",x"C9",x"2C",x"D0",x"1E",x"20", -- 0x06E8
    x"2C",x"88",x"20",x"97",x"8A",x"C9",x"59",x"D0", -- 0x06F0
    x"14",x"F0",x"CD",x"C9",x"2C",x"D0",x"0E",x"20", -- 0x06F8
    x"97",x"8A",x"C9",x"58",x"D0",x"07",x"20",x"97", -- 0x0700
    x"8A",x"C9",x"29",x"F0",x"BB",x"00",x"03",x"49", -- 0x0708
    x"6E",x"64",x"65",x"78",x"00",x"C6",x"0A",x"20", -- 0x0710
    x"21",x"88",x"20",x"97",x"8A",x"C9",x"2C",x"D0", -- 0x0718
    x"14",x"20",x"2C",x"88",x"20",x"97",x"8A",x"C9", -- 0x0720
    x"58",x"F0",x"0A",x"C9",x"59",x"D0",x"DE",x"20", -- 0x0728
    x"2F",x"88",x"4C",x"9A",x"87",x"20",x"32",x"88", -- 0x0730
    x"A5",x"2B",x"D0",x"F3",x"4C",x"A8",x"86",x"E0", -- 0x0738
    x"2F",x"B0",x"2B",x"E0",x"2D",x"B0",x"09",x"20", -- 0x0740
    x"97",x"8A",x"C9",x"41",x"F0",x"19",x"C6",x"0A", -- 0x0748
    x"20",x"21",x"88",x"20",x"97",x"8A",x"C9",x"2C", -- 0x0750
    x"D0",x"DE",x"20",x"2C",x"88",x"20",x"97",x"8A", -- 0x0758
    x"C9",x"58",x"F0",x"D4",x"4C",x"0D",x"87",x"20", -- 0x0760
    x"32",x"88",x"A0",x"01",x"D0",x"2E",x"E0",x"32", -- 0x0768
    x"B0",x"16",x"E0",x"31",x"F0",x"0C",x"20",x"97", -- 0x0770
    x"8A",x"C9",x"23",x"D0",x"03",x"4C",x"C5",x"86", -- 0x0778
    x"C6",x"0A",x"20",x"21",x"88",x"4C",x"35",x"87", -- 0x0780
    x"E0",x"33",x"F0",x"0B",x"B0",x"24",x"20",x"97", -- 0x0788
    x"8A",x"C9",x"28",x"F0",x"0A",x"C6",x"0A",x"20", -- 0x0790
    x"21",x"88",x"A0",x"03",x"4C",x"2B",x"86",x"20", -- 0x0798
    x"2C",x"88",x"20",x"2C",x"88",x"20",x"21",x"88", -- 0x07A0
    x"20",x"97",x"8A",x"C9",x"29",x"F0",x"EB",x"4C", -- 0x07A8
    x"0D",x"87",x"E0",x"39",x"B0",x"5D",x"A5",x"3D", -- 0x07B0
    x"49",x"01",x"29",x"1F",x"48",x"E0",x"37",x"B0", -- 0x07B8
    x"2F",x"20",x"97",x"8A",x"C9",x"23",x"D0",x"04", -- 0x07C0
    x"68",x"4C",x"C5",x"86",x"C6",x"0A",x"20",x"21", -- 0x07C8
    x"88",x"68",x"85",x"37",x"20",x"97",x"8A",x"C9", -- 0x07D0
    x"2C",x"F0",x"03",x"4C",x"35",x"87",x"20",x"97", -- 0x07D8
    x"8A",x"29",x"1F",x"C5",x"37",x"D0",x"06",x"20", -- 0x07E0
    x"2C",x"88",x"4C",x"35",x"87",x"4C",x"0D",x"87", -- 0x07E8
    x"20",x"21",x"88",x"68",x"85",x"37",x"20",x"97", -- 0x07F0
    x"8A",x"C9",x"2C",x"D0",x"13",x"20",x"97",x"8A", -- 0x07F8
    x"29",x"1F",x"C5",x"37",x"D0",x"E7",x"20",x"2C", -- 0x0800
    x"88",x"A5",x"2B",x"F0",x"03",x"4C",x"CC",x"86", -- 0x0808
    x"4C",x"38",x"87",x"D0",x"25",x"20",x"21",x"88", -- 0x0810
    x"A5",x"2A",x"85",x"28",x"A0",x"00",x"4C",x"2B", -- 0x0818
    x"86",x"20",x"1D",x"9B",x"20",x"F0",x"92",x"A4", -- 0x0820
    x"1B",x"84",x"0A",x"60",x"20",x"2F",x"88",x"20", -- 0x0828
    x"32",x"88",x"A5",x"29",x"18",x"69",x"04",x"85", -- 0x0830
    x"29",x"60",x"A2",x"01",x"A4",x"0A",x"E6",x"0A", -- 0x0838
    x"B1",x"0B",x"C9",x"42",x"F0",x"12",x"E8",x"C9", -- 0x0840
    x"57",x"F0",x"0D",x"A2",x"04",x"C9",x"44",x"F0", -- 0x0848
    x"07",x"C9",x"53",x"F0",x"15",x"4C",x"2A",x"98", -- 0x0850
    x"8A",x"48",x"20",x"21",x"88",x"A2",x"29",x"20", -- 0x0858
    x"44",x"BE",x"68",x"A8",x"4C",x"2B",x"86",x"4C", -- 0x0860
    x"0E",x"8C",x"A5",x"28",x"48",x"20",x"1D",x"9B", -- 0x0868
    x"D0",x"F5",x"68",x"85",x"28",x"20",x"27",x"88", -- 0x0870
    x"A0",x"FF",x"D0",x"E8",x"48",x"18",x"98",x"65", -- 0x0878
    x"37",x"85",x"39",x"A0",x"00",x"98",x"65",x"38", -- 0x0880
    x"85",x"3A",x"68",x"91",x"37",x"C8",x"B1",x"39", -- 0x0888
    x"91",x"37",x"C9",x"0D",x"D0",x"F7",x"60",x"29", -- 0x0890
    x"0F",x"85",x"3D",x"84",x"3E",x"C8",x"B1",x"37", -- 0x0898
    x"C9",x"3A",x"B0",x"36",x"C9",x"30",x"90",x"32", -- 0x08A0
    x"29",x"0F",x"48",x"A6",x"3E",x"A5",x"3D",x"0A", -- 0x08A8
    x"26",x"3E",x"30",x"21",x"0A",x"26",x"3E",x"30", -- 0x08B0
    x"1C",x"65",x"3D",x"85",x"3D",x"8A",x"65",x"3E", -- 0x08B8
    x"06",x"3D",x"2A",x"30",x"10",x"B0",x"0E",x"85", -- 0x08C0
    x"3E",x"68",x"65",x"3D",x"85",x"3D",x"90",x"CD", -- 0x08C8
    x"E6",x"3E",x"10",x"C9",x"48",x"68",x"A0",x"00", -- 0x08D0
    x"38",x"60",x"88",x"A9",x"8D",x"20",x"7C",x"88", -- 0x08D8
    x"A5",x"37",x"69",x"02",x"85",x"39",x"A5",x"38", -- 0x08E0
    x"69",x"00",x"85",x"3A",x"B1",x"37",x"91",x"39", -- 0x08E8
    x"88",x"D0",x"F9",x"A0",x"03",x"A5",x"3E",x"09", -- 0x08F0
    x"40",x"91",x"37",x"88",x"A5",x"3D",x"29",x"3F", -- 0x08F8
    x"09",x"40",x"91",x"37",x"88",x"A5",x"3D",x"29", -- 0x0900
    x"C0",x"85",x"3D",x"A5",x"3E",x"29",x"C0",x"4A", -- 0x0908
    x"4A",x"05",x"3D",x"4A",x"4A",x"49",x"54",x"91", -- 0x0910
    x"37",x"20",x"44",x"89",x"20",x"44",x"89",x"20", -- 0x0918
    x"44",x"89",x"A0",x"00",x"18",x"60",x"C9",x"7B", -- 0x0920
    x"B0",x"FA",x"C9",x"5F",x"B0",x"0E",x"C9",x"5B", -- 0x0928
    x"B0",x"F2",x"C9",x"41",x"B0",x"06",x"C9",x"3A", -- 0x0930
    x"B0",x"EA",x"C9",x"30",x"60",x"C9",x"2E",x"D0", -- 0x0938
    x"F5",x"60",x"B1",x"37",x"E6",x"37",x"D0",x"02", -- 0x0940
    x"E6",x"38",x"60",x"20",x"44",x"89",x"B1",x"37", -- 0x0948
    x"60",x"A0",x"00",x"84",x"3B",x"84",x"3C",x"B1", -- 0x0950
    x"37",x"C9",x"0D",x"F0",x"ED",x"C9",x"20",x"D0", -- 0x0958
    x"05",x"20",x"44",x"89",x"D0",x"F1",x"C9",x"26", -- 0x0960
    x"D0",x"12",x"20",x"4B",x"89",x"20",x"36",x"89", -- 0x0968
    x"B0",x"F8",x"C9",x"41",x"90",x"E1",x"C9",x"47", -- 0x0970
    x"90",x"F0",x"B0",x"DB",x"C9",x"22",x"D0",x"0C", -- 0x0978
    x"20",x"4B",x"89",x"C9",x"22",x"F0",x"DA",x"C9", -- 0x0980
    x"0D",x"D0",x"F5",x"60",x"C9",x"3A",x"D0",x"06", -- 0x0988
    x"84",x"3B",x"84",x"3C",x"F0",x"CB",x"C9",x"2C", -- 0x0990
    x"F0",x"C7",x"C9",x"2A",x"D0",x"05",x"A5",x"3B", -- 0x0998
    x"D0",x"41",x"60",x"C9",x"2E",x"F0",x"0E",x"20", -- 0x09A0
    x"36",x"89",x"90",x"33",x"A6",x"3C",x"F0",x"05", -- 0x09A8
    x"20",x"97",x"88",x"90",x"34",x"B1",x"37",x"20", -- 0x09B0
    x"3D",x"89",x"90",x"06",x"20",x"44",x"89",x"4C", -- 0x09B8
    x"B5",x"89",x"A2",x"FF",x"86",x"3B",x"84",x"3C", -- 0x09C0
    x"4C",x"57",x"89",x"20",x"26",x"89",x"90",x"13", -- 0x09C8
    x"A0",x"00",x"B1",x"37",x"20",x"26",x"89",x"90", -- 0x09D0
    x"E9",x"20",x"44",x"89",x"4C",x"D2",x"89",x"C9", -- 0x09D8
    x"41",x"B0",x"09",x"A2",x"FF",x"86",x"3B",x"84", -- 0x09E0
    x"3C",x"4C",x"61",x"89",x"C9",x"58",x"B0",x"DB", -- 0x09E8
    x"A2",x"71",x"86",x"39",x"A2",x"80",x"86",x"3A", -- 0x09F0
    x"D1",x"39",x"90",x"D6",x"D0",x"0F",x"C8",x"B1", -- 0x09F8
    x"39",x"30",x"34",x"D1",x"37",x"F0",x"F7",x"B1", -- 0x0A00
    x"37",x"C9",x"2E",x"F0",x"0B",x"C8",x"B1",x"39", -- 0x0A08
    x"10",x"FB",x"C9",x"FE",x"D0",x"0F",x"B0",x"B8", -- 0x0A10
    x"C8",x"B1",x"39",x"30",x"1A",x"E6",x"39",x"D0", -- 0x0A18
    x"F8",x"E6",x"3A",x"D0",x"F4",x"38",x"C8",x"98", -- 0x0A20
    x"65",x"39",x"85",x"39",x"90",x"02",x"E6",x"3A", -- 0x0A28
    x"A0",x"00",x"B1",x"37",x"4C",x"F8",x"89",x"AA", -- 0x0A30
    x"C8",x"B1",x"39",x"85",x"3D",x"88",x"4A",x"90", -- 0x0A38
    x"07",x"B1",x"37",x"20",x"26",x"89",x"B0",x"88", -- 0x0A40
    x"8A",x"24",x"3D",x"50",x"07",x"A6",x"3B",x"D0", -- 0x0A48
    x"03",x"18",x"69",x"40",x"88",x"20",x"7C",x"88", -- 0x0A50
    x"A0",x"00",x"A2",x"FF",x"A5",x"3D",x"4A",x"4A", -- 0x0A58
    x"90",x"04",x"86",x"3B",x"84",x"3C",x"4A",x"90", -- 0x0A60
    x"04",x"84",x"3B",x"84",x"3C",x"4A",x"90",x"11", -- 0x0A68
    x"48",x"C8",x"B1",x"37",x"20",x"26",x"89",x"90", -- 0x0A70
    x"06",x"20",x"44",x"89",x"4C",x"72",x"8A",x"88", -- 0x0A78
    x"68",x"4A",x"90",x"02",x"86",x"3C",x"4A",x"B0", -- 0x0A80
    x"0D",x"4C",x"61",x"89",x"A4",x"1B",x"E6",x"1B", -- 0x0A88
    x"B1",x"19",x"C9",x"20",x"F0",x"F6",x"60",x"A4", -- 0x0A90
    x"0A",x"E6",x"0A",x"B1",x"0B",x"C9",x"20",x"F0", -- 0x0A98
    x"F6",x"60",x"00",x"05",x"4D",x"69",x"73",x"73", -- 0x0AA0
    x"69",x"6E",x"67",x"20",x"2C",x"00",x"20",x"8C", -- 0x0AA8
    x"8A",x"C9",x"2C",x"D0",x"ED",x"60",x"20",x"57", -- 0x0AB0
    x"98",x"A5",x"18",x"85",x"38",x"A9",x"00",x"85", -- 0x0AB8
    x"37",x"91",x"37",x"20",x"6F",x"BE",x"D0",x"2B", -- 0x0AC0
    x"20",x"57",x"98",x"20",x"6F",x"BE",x"D0",x"26", -- 0x0AC8
    x"20",x"57",x"98",x"00",x"00",x"53",x"54",x"4F", -- 0x0AD0
    x"50",x"00",x"20",x"57",x"98",x"A9",x"0D",x"A4", -- 0x0AD8
    x"18",x"84",x"13",x"A0",x"00",x"84",x"12",x"84", -- 0x0AE0
    x"20",x"91",x"12",x"A9",x"FF",x"C8",x"91",x"12", -- 0x0AE8
    x"C8",x"84",x"12",x"20",x"20",x"BD",x"A0",x"07", -- 0x0AF0
    x"84",x"0C",x"A0",x"00",x"84",x"0B",x"A9",x"33", -- 0x0AF8
    x"85",x"16",x"A9",x"B4",x"85",x"17",x"A9",x"3E", -- 0x0B00
    x"20",x"02",x"BC",x"A9",x"33",x"85",x"16",x"A9", -- 0x0B08
    x"B4",x"85",x"17",x"A2",x"FF",x"86",x"28",x"86", -- 0x0B10
    x"3C",x"9A",x"20",x"3A",x"BD",x"A8",x"A5",x"0B", -- 0x0B18
    x"85",x"37",x"A5",x"0C",x"85",x"38",x"84",x"3B", -- 0x0B20
    x"84",x"0A",x"20",x"57",x"89",x"20",x"DF",x"97", -- 0x0B28
    x"90",x"06",x"20",x"8D",x"BC",x"4C",x"F3",x"8A", -- 0x0B30
    x"20",x"97",x"8A",x"C9",x"C6",x"B0",x"72",x"90", -- 0x0B38
    x"7E",x"4C",x"F6",x"8A",x"4C",x"04",x"85",x"BA", -- 0x0B40
    x"E0",x"FC",x"B0",x"0D",x"AD",x"FF",x"01",x"C9", -- 0x0B48
    x"A4",x"D0",x"06",x"20",x"1D",x"9B",x"4C",x"4C", -- 0x0B50
    x"98",x"00",x"07",x"4E",x"6F",x"20",x"A4",x"00", -- 0x0B58
    x"A4",x"0A",x"88",x"B1",x"0B",x"C9",x"3D",x"F0", -- 0x0B60
    x"DE",x"C9",x"2A",x"F0",x"06",x"C9",x"5B",x"F0", -- 0x0B68
    x"D3",x"D0",x"23",x"20",x"6D",x"98",x"A6",x"0B", -- 0x0B70
    x"A4",x"0C",x"20",x"F7",x"FF",x"A9",x"0D",x"A4", -- 0x0B78
    x"0A",x"88",x"C8",x"D1",x"0B",x"D0",x"FB",x"C9", -- 0x0B80
    x"8B",x"F0",x"F2",x"A5",x"0C",x"C9",x"07",x"F0", -- 0x0B88
    x"B0",x"20",x"90",x"98",x"D0",x"0D",x"C6",x"0A", -- 0x0B90
    x"20",x"57",x"98",x"A0",x"00",x"B1",x"0B",x"C9", -- 0x0B98
    x"3A",x"D0",x"E4",x"A4",x"0A",x"E6",x"0A",x"B1", -- 0x0BA0
    x"0B",x"C9",x"20",x"F0",x"F6",x"C9",x"CF",x"90", -- 0x0BA8
    x"0E",x"AA",x"BD",x"DF",x"82",x"85",x"37",x"BD", -- 0x0BB0
    x"51",x"83",x"85",x"38",x"6C",x"37",x"00",x"A6", -- 0x0BB8
    x"0B",x"86",x"19",x"A6",x"0C",x"86",x"1A",x"84", -- 0x0BC0
    x"1B",x"20",x"DD",x"95",x"D0",x"1B",x"B0",x"90", -- 0x0BC8
    x"86",x"1B",x"20",x"41",x"98",x"20",x"FC",x"94", -- 0x0BD0
    x"A2",x"05",x"E4",x"2C",x"D0",x"01",x"E8",x"20", -- 0x0BD8
    x"31",x"95",x"C6",x"0A",x"20",x"82",x"95",x"F0", -- 0x0BE0
    x"22",x"90",x"10",x"20",x"94",x"BD",x"20",x"13", -- 0x0BE8
    x"98",x"A5",x"27",x"D0",x"19",x"20",x"1E",x"8C", -- 0x0BF0
    x"4C",x"9B",x"8B",x"20",x"94",x"BD",x"20",x"13", -- 0x0BF8
    x"98",x"A5",x"27",x"F0",x"09",x"20",x"B4",x"B4", -- 0x0C00
    x"4C",x"9B",x"8B",x"4C",x"2A",x"98",x"00",x"06", -- 0x0C08
    x"54",x"79",x"70",x"65",x"20",x"6D",x"69",x"73", -- 0x0C10
    x"6D",x"61",x"74",x"63",x"68",x"00",x"20",x"EA", -- 0x0C18
    x"BD",x"A5",x"2C",x"C9",x"80",x"F0",x"7B",x"A0", -- 0x0C20
    x"02",x"B1",x"2A",x"C5",x"36",x"B0",x"55",x"A5", -- 0x0C28
    x"02",x"85",x"2C",x"A5",x"03",x"85",x"2D",x"A5", -- 0x0C30
    x"36",x"C9",x"08",x"90",x"06",x"69",x"07",x"90", -- 0x0C38
    x"02",x"A9",x"FF",x"18",x"48",x"AA",x"B1",x"2A", -- 0x0C40
    x"A0",x"00",x"71",x"2A",x"45",x"02",x"D0",x"0F", -- 0x0C48
    x"C8",x"71",x"2A",x"45",x"03",x"D0",x"08",x"85", -- 0x0C50
    x"2D",x"8A",x"C8",x"38",x"F1",x"2A",x"AA",x"8A", -- 0x0C58
    x"18",x"65",x"02",x"A8",x"A5",x"03",x"69",x"00", -- 0x0C60
    x"C4",x"04",x"AA",x"E5",x"05",x"B0",x"48",x"84", -- 0x0C68
    x"02",x"86",x"03",x"68",x"A0",x"02",x"91",x"2A", -- 0x0C70
    x"88",x"A5",x"2D",x"F0",x"07",x"91",x"2A",x"88", -- 0x0C78
    x"A5",x"2C",x"91",x"2A",x"A0",x"03",x"A5",x"36", -- 0x0C80
    x"91",x"2A",x"F0",x"15",x"88",x"88",x"B1",x"2A", -- 0x0C88
    x"85",x"2D",x"88",x"B1",x"2A",x"85",x"2C",x"B9", -- 0x0C90
    x"00",x"06",x"91",x"2C",x"C8",x"C4",x"36",x"D0", -- 0x0C98
    x"F6",x"60",x"20",x"BA",x"BE",x"C0",x"00",x"F0", -- 0x0CA0
    x"0B",x"B9",x"00",x"06",x"91",x"2A",x"88",x"D0", -- 0x0CA8
    x"F8",x"AD",x"00",x"06",x"91",x"2A",x"60",x"00", -- 0x0CB0
    x"00",x"4E",x"6F",x"20",x"72",x"6F",x"6F",x"6D", -- 0x0CB8
    x"00",x"A5",x"39",x"C9",x"80",x"F0",x"27",x"90", -- 0x0CC0
    x"3A",x"A0",x"00",x"B1",x"04",x"AA",x"F0",x"15", -- 0x0CC8
    x"B1",x"37",x"E9",x"01",x"85",x"39",x"C8",x"B1", -- 0x0CD0
    x"37",x"E9",x"00",x"85",x"3A",x"B1",x"04",x"91", -- 0x0CD8
    x"39",x"C8",x"CA",x"D0",x"F8",x"A1",x"04",x"A0", -- 0x0CE0
    x"03",x"91",x"37",x"4C",x"DC",x"BD",x"A0",x"00", -- 0x0CE8
    x"B1",x"04",x"AA",x"F0",x"0A",x"C8",x"B1",x"04", -- 0x0CF0
    x"88",x"91",x"37",x"C8",x"CA",x"D0",x"F6",x"A9", -- 0x0CF8
    x"0D",x"D0",x"E6",x"A0",x"00",x"B1",x"04",x"91", -- 0x0D00
    x"37",x"C8",x"C4",x"39",x"B0",x"18",x"B1",x"04", -- 0x0D08
    x"91",x"37",x"C8",x"B1",x"04",x"91",x"37",x"C8", -- 0x0D10
    x"B1",x"04",x"91",x"37",x"C8",x"C4",x"39",x"B0", -- 0x0D18
    x"05",x"B1",x"04",x"91",x"37",x"C8",x"98",x"18", -- 0x0D20
    x"4C",x"E1",x"BD",x"C6",x"0A",x"20",x"A9",x"BF", -- 0x0D28
    x"98",x"48",x"20",x"8C",x"8A",x"C9",x"2C",x"D0", -- 0x0D30
    x"3E",x"20",x"29",x"9B",x"20",x"85",x"A3",x"68", -- 0x0D38
    x"A8",x"A5",x"27",x"20",x"D4",x"FF",x"AA",x"F0", -- 0x0D40
    x"1B",x"30",x"0C",x"A2",x"03",x"B5",x"2A",x"20", -- 0x0D48
    x"D4",x"FF",x"CA",x"10",x"F8",x"30",x"D9",x"A2", -- 0x0D50
    x"04",x"BD",x"6C",x"04",x"20",x"D4",x"FF",x"CA", -- 0x0D58
    x"10",x"F7",x"30",x"CC",x"A5",x"36",x"20",x"D4", -- 0x0D60
    x"FF",x"AA",x"F0",x"C4",x"BD",x"FF",x"05",x"20", -- 0x0D68
    x"D4",x"FF",x"CA",x"D0",x"F7",x"F0",x"B9",x"68", -- 0x0D70
    x"84",x"0A",x"4C",x"98",x"8B",x"20",x"25",x"BC", -- 0x0D78
    x"4C",x"96",x"8B",x"A9",x"00",x"85",x"14",x"85", -- 0x0D80
    x"15",x"20",x"97",x"8A",x"C9",x"3A",x"F0",x"F0", -- 0x0D88
    x"C9",x"0D",x"F0",x"EC",x"C9",x"8B",x"F0",x"E8", -- 0x0D90
    x"D0",x"38",x"20",x"97",x"8A",x"C9",x"23",x"F0", -- 0x0D98
    x"8A",x"C6",x"0A",x"4C",x"BB",x"8D",x"AD",x"00", -- 0x0DA0
    x"04",x"F0",x"10",x"A5",x"1E",x"F0",x"0C",x"ED", -- 0x0DA8
    x"00",x"04",x"B0",x"F9",x"A8",x"20",x"65",x"B5", -- 0x0DB0
    x"C8",x"D0",x"FA",x"18",x"AD",x"00",x"04",x"85", -- 0x0DB8
    x"14",x"66",x"15",x"20",x"97",x"8A",x"C9",x"3A", -- 0x0DC0
    x"F0",x"B3",x"C9",x"0D",x"F0",x"AF",x"C9",x"8B", -- 0x0DC8
    x"F0",x"AB",x"C9",x"7E",x"F0",x"EB",x"C9",x"2C", -- 0x0DD0
    x"F0",x"CC",x"C9",x"3B",x"F0",x"A5",x"20",x"70", -- 0x0DD8
    x"8E",x"90",x"E0",x"A5",x"14",x"48",x"A5",x"15", -- 0x0DE0
    x"48",x"C6",x"1B",x"20",x"29",x"9B",x"68",x"85", -- 0x0DE8
    x"15",x"68",x"85",x"14",x"A5",x"1B",x"85",x"0A", -- 0x0DF0
    x"98",x"F0",x"13",x"20",x"DF",x"9E",x"A5",x"14", -- 0x0DF8
    x"38",x"E5",x"36",x"90",x"09",x"F0",x"07",x"A8", -- 0x0E00
    x"20",x"65",x"B5",x"88",x"D0",x"FA",x"A5",x"36", -- 0x0E08
    x"F0",x"B1",x"A0",x"00",x"B9",x"00",x"06",x"20", -- 0x0E10
    x"58",x"B5",x"C8",x"C4",x"36",x"D0",x"F5",x"F0", -- 0x0E18
    x"A2",x"4C",x"A2",x"8A",x"C9",x"2C",x"D0",x"F9", -- 0x0E20
    x"A5",x"2A",x"48",x"20",x"56",x"AE",x"20",x"F0", -- 0x0E28
    x"92",x"A9",x"1F",x"20",x"EE",x"FF",x"68",x"20", -- 0x0E30
    x"EE",x"FF",x"20",x"56",x"94",x"4C",x"6A",x"8E", -- 0x0E38
    x"20",x"DD",x"92",x"20",x"8C",x"8A",x"C9",x"29", -- 0x0E40
    x"D0",x"DA",x"A5",x"2A",x"E5",x"1E",x"F0",x"1A", -- 0x0E48
    x"A8",x"B0",x"0C",x"20",x"25",x"BC",x"F0",x"03", -- 0x0E50
    x"20",x"E3",x"92",x"A4",x"2A",x"F0",x"0B",x"20", -- 0x0E58
    x"65",x"B5",x"88",x"D0",x"FA",x"F0",x"03",x"20", -- 0x0E60
    x"25",x"BC",x"18",x"A4",x"1B",x"84",x"0A",x"60", -- 0x0E68
    x"A6",x"0B",x"86",x"19",x"A6",x"0C",x"86",x"1A", -- 0x0E70
    x"A6",x"0A",x"86",x"1B",x"C9",x"27",x"F0",x"E7", -- 0x0E78
    x"C9",x"8A",x"F0",x"BC",x"C9",x"89",x"F0",x"D0", -- 0x0E80
    x"38",x"60",x"20",x"97",x"8A",x"20",x"70",x"8E", -- 0x0E88
    x"90",x"F7",x"C9",x"22",x"F0",x"11",x"38",x"60", -- 0x0E90
    x"00",x"09",x"4D",x"69",x"73",x"73",x"69",x"6E", -- 0x0E98
    x"67",x"20",x"22",x"00",x"20",x"58",x"B5",x"C8", -- 0x0EA0
    x"B1",x"19",x"C9",x"0D",x"F0",x"EA",x"C9",x"22", -- 0x0EA8
    x"D0",x"F2",x"C8",x"84",x"1B",x"B1",x"19",x"C9", -- 0x0EB0
    x"22",x"D0",x"AF",x"F0",x"E7",x"20",x"57",x"98", -- 0x0EB8
    x"A9",x"10",x"D0",x"08",x"20",x"57",x"98",x"20", -- 0x0EC0
    x"28",x"BC",x"A9",x"0C",x"20",x"EE",x"FF",x"4C", -- 0x0EC8
    x"9B",x"8B",x"20",x"1D",x"9B",x"20",x"EE",x"92", -- 0x0ED0
    x"20",x"94",x"BD",x"A0",x"00",x"8C",x"00",x"06", -- 0x0ED8
    x"8C",x"FF",x"06",x"20",x"8C",x"8A",x"C9",x"2C", -- 0x0EE0
    x"D0",x"22",x"A4",x"1B",x"20",x"D5",x"95",x"F0", -- 0x0EE8
    x"2A",x"AC",x"FF",x"06",x"C8",x"A5",x"2A",x"99", -- 0x0EF0
    x"00",x"06",x"C8",x"A5",x"2B",x"99",x"00",x"06", -- 0x0EF8
    x"C8",x"A5",x"2C",x"99",x"00",x"06",x"EE",x"00", -- 0x0F00
    x"06",x"4C",x"E0",x"8E",x"C6",x"1B",x"20",x"52", -- 0x0F08
    x"98",x"20",x"EA",x"BD",x"20",x"1E",x"8F",x"D8", -- 0x0F10
    x"4C",x"9B",x"8B",x"4C",x"43",x"AE",x"AD",x"0C", -- 0x0F18
    x"04",x"4A",x"AD",x"04",x"04",x"AE",x"60",x"04", -- 0x0F20
    x"AC",x"64",x"04",x"6C",x"2A",x"00",x"4C",x"2A", -- 0x0F28
    x"98",x"20",x"DF",x"97",x"90",x"F8",x"20",x"94", -- 0x0F30
    x"BD",x"20",x"97",x"8A",x"C9",x"2C",x"D0",x"EE", -- 0x0F38
    x"20",x"DF",x"97",x"90",x"E9",x"20",x"57",x"98", -- 0x0F40
    x"A5",x"2A",x"85",x"39",x"A5",x"2B",x"85",x"3A", -- 0x0F48
    x"20",x"EA",x"BD",x"20",x"2D",x"BC",x"20",x"7B", -- 0x0F50
    x"98",x"20",x"22",x"92",x"A5",x"39",x"C5",x"2A", -- 0x0F58
    x"A5",x"3A",x"E5",x"2B",x"B0",x"ED",x"4C",x"F3", -- 0x0F60
    x"8A",x"A9",x"0A",x"20",x"D8",x"AE",x"20",x"DF", -- 0x0F68
    x"97",x"20",x"94",x"BD",x"A9",x"0A",x"20",x"D8", -- 0x0F70
    x"AE",x"20",x"97",x"8A",x"C9",x"2C",x"D0",x"0D", -- 0x0F78
    x"20",x"DF",x"97",x"A5",x"2B",x"D0",x"58",x"A5", -- 0x0F80
    x"2A",x"F0",x"54",x"E6",x"0A",x"C6",x"0A",x"4C", -- 0x0F88
    x"57",x"98",x"A5",x"12",x"85",x"3B",x"A5",x"13", -- 0x0F90
    x"85",x"3C",x"A5",x"18",x"85",x"38",x"A9",x"01", -- 0x0F98
    x"85",x"37",x"60",x"20",x"69",x"8F",x"A2",x"39", -- 0x0FA0
    x"20",x"0D",x"BE",x"20",x"6F",x"BE",x"20",x"92", -- 0x0FA8
    x"8F",x"A0",x"00",x"B1",x"37",x"30",x"30",x"91", -- 0x0FB0
    x"3B",x"C8",x"B1",x"37",x"91",x"3B",x"38",x"98", -- 0x0FB8
    x"65",x"3B",x"85",x"3B",x"AA",x"A5",x"3C",x"69", -- 0x0FC0
    x"00",x"85",x"3C",x"E4",x"06",x"E5",x"07",x"B0", -- 0x0FC8
    x"05",x"20",x"9F",x"90",x"90",x"DB",x"00",x"00", -- 0x0FD0
    x"CC",x"20",x"73",x"70",x"61",x"63",x"65",x"00", -- 0x0FD8
    x"00",x"53",x"69",x"6C",x"6C",x"79",x"00",x"20", -- 0x0FE0
    x"9A",x"8F",x"A0",x"00",x"B1",x"37",x"30",x"1D", -- 0x0FE8
    x"A5",x"3A",x"91",x"37",x"A5",x"39",x"C8",x"91", -- 0x0FF0
    x"37",x"18",x"A5",x"2A",x"65",x"39",x"85",x"39", -- 0x0FF8
    x"A9",x"00",x"65",x"3A",x"29",x"7F",x"85",x"3A", -- 0x1000
    x"20",x"9F",x"90",x"90",x"DD",x"A5",x"18",x"85", -- 0x1008
    x"0C",x"A0",x"00",x"84",x"0B",x"C8",x"B1",x"0B", -- 0x1010
    x"30",x"20",x"A0",x"04",x"B1",x"0B",x"C9",x"8D", -- 0x1018
    x"F0",x"1B",x"C8",x"C9",x"0D",x"D0",x"F5",x"B1", -- 0x1020
    x"0B",x"30",x"0F",x"A0",x"03",x"B1",x"0B",x"18", -- 0x1028
    x"65",x"0B",x"85",x"0B",x"90",x"E4",x"E6",x"0C", -- 0x1030
    x"B0",x"E0",x"4C",x"F3",x"8A",x"20",x"EB",x"97", -- 0x1038
    x"20",x"92",x"8F",x"A0",x"00",x"B1",x"37",x"30", -- 0x1040
    x"37",x"B1",x"3B",x"C8",x"C5",x"2B",x"D0",x"21", -- 0x1048
    x"B1",x"3B",x"C5",x"2A",x"D0",x"1B",x"B1",x"37", -- 0x1050
    x"85",x"3D",x"88",x"B1",x"37",x"85",x"3E",x"A4", -- 0x1058
    x"0A",x"88",x"A5",x"0B",x"85",x"37",x"A5",x"0C", -- 0x1060
    x"85",x"38",x"20",x"F5",x"88",x"A4",x"0A",x"D0", -- 0x1068
    x"AB",x"20",x"9F",x"90",x"A5",x"3B",x"69",x"02", -- 0x1070
    x"85",x"3B",x"90",x"C7",x"E6",x"3C",x"B0",x"C3", -- 0x1078
    x"20",x"CF",x"BF",x"46",x"61",x"69",x"6C",x"65", -- 0x1080
    x"64",x"20",x"61",x"74",x"20",x"C8",x"B1",x"0B", -- 0x1088
    x"85",x"2B",x"C8",x"B1",x"0B",x"85",x"2A",x"20", -- 0x1090
    x"1F",x"99",x"20",x"25",x"BC",x"F0",x"CE",x"C8", -- 0x1098
    x"B1",x"37",x"65",x"37",x"85",x"37",x"90",x"03", -- 0x10A0
    x"E6",x"38",x"18",x"60",x"20",x"69",x"8F",x"A5", -- 0x10A8
    x"2A",x"48",x"20",x"EA",x"BD",x"20",x"94",x"BD", -- 0x10B0
    x"20",x"23",x"99",x"A9",x"20",x"20",x"02",x"BC", -- 0x10B8
    x"20",x"EA",x"BD",x"20",x"51",x"89",x"20",x"8D", -- 0x10C0
    x"BC",x"20",x"20",x"BD",x"68",x"48",x"18",x"65", -- 0x10C8
    x"2A",x"85",x"2A",x"90",x"E0",x"E6",x"2B",x"10", -- 0x10D0
    x"DC",x"4C",x"F3",x"8A",x"4C",x"18",x"92",x"C6", -- 0x10D8
    x"0A",x"20",x"82",x"95",x"F0",x"41",x"B0",x"3F", -- 0x10E0
    x"20",x"94",x"BD",x"20",x"DD",x"92",x"20",x"22", -- 0x10E8
    x"92",x"A5",x"2D",x"05",x"2C",x"D0",x"30",x"18", -- 0x10F0
    x"A5",x"2A",x"65",x"02",x"A8",x"A5",x"2B",x"65", -- 0x10F8
    x"03",x"AA",x"C4",x"04",x"E5",x"05",x"B0",x"D4", -- 0x1100
    x"A5",x"02",x"85",x"2A",x"A5",x"03",x"85",x"2B", -- 0x1108
    x"84",x"02",x"86",x"03",x"A9",x"00",x"85",x"2C", -- 0x1110
    x"85",x"2D",x"A9",x"40",x"85",x"27",x"20",x"B4", -- 0x1118
    x"B4",x"20",x"27",x"88",x"4C",x"0B",x"92",x"00", -- 0x1120
    x"0A",x"42",x"61",x"64",x"20",x"DE",x"00",x"20", -- 0x1128
    x"97",x"8A",x"98",x"18",x"65",x"0B",x"A6",x"0C", -- 0x1130
    x"90",x"02",x"E8",x"18",x"E9",x"00",x"85",x"37", -- 0x1138
    x"8A",x"E9",x"00",x"85",x"38",x"A2",x"05",x"86", -- 0x1140
    x"3F",x"A6",x"0A",x"20",x"59",x"95",x"C0",x"01", -- 0x1148
    x"F0",x"D5",x"C9",x"28",x"F0",x"15",x"C9",x"24", -- 0x1150
    x"F0",x"04",x"C9",x"25",x"D0",x"0A",x"C6",x"3F", -- 0x1158
    x"C8",x"E8",x"B1",x"37",x"C9",x"28",x"F0",x"03", -- 0x1160
    x"4C",x"DF",x"90",x"84",x"39",x"86",x"0A",x"20", -- 0x1168
    x"69",x"94",x"D0",x"B3",x"20",x"FC",x"94",x"A2", -- 0x1170
    x"01",x"20",x"31",x"95",x"A5",x"3F",x"48",x"A9", -- 0x1178
    x"01",x"48",x"20",x"D8",x"AE",x"20",x"94",x"BD", -- 0x1180
    x"20",x"21",x"88",x"A5",x"2B",x"29",x"C0",x"05", -- 0x1188
    x"2C",x"05",x"2D",x"D0",x"92",x"20",x"22",x"92", -- 0x1190
    x"68",x"A8",x"A5",x"2A",x"91",x"02",x"C8",x"A5", -- 0x1198
    x"2B",x"91",x"02",x"C8",x"98",x"48",x"20",x"31", -- 0x11A0
    x"92",x"20",x"97",x"8A",x"C9",x"2C",x"F0",x"D5", -- 0x11A8
    x"C9",x"29",x"F0",x"03",x"4C",x"27",x"91",x"68", -- 0x11B0
    x"85",x"15",x"68",x"85",x"3F",x"A9",x"00",x"85", -- 0x11B8
    x"40",x"20",x"36",x"92",x"A0",x"00",x"A5",x"15", -- 0x11C0
    x"91",x"02",x"65",x"2A",x"85",x"2A",x"90",x"02", -- 0x11C8
    x"E6",x"2B",x"A5",x"03",x"85",x"38",x"A5",x"02", -- 0x11D0
    x"85",x"37",x"18",x"65",x"2A",x"A8",x"A5",x"2B", -- 0x11D8
    x"65",x"03",x"B0",x"34",x"AA",x"C4",x"04",x"E5", -- 0x11E0
    x"05",x"B0",x"2D",x"84",x"02",x"86",x"03",x"A5", -- 0x11E8
    x"37",x"65",x"15",x"A8",x"A9",x"00",x"85",x"37", -- 0x11F0
    x"90",x"02",x"E6",x"38",x"91",x"37",x"C8",x"D0", -- 0x11F8
    x"02",x"E6",x"38",x"C4",x"02",x"D0",x"F5",x"E4", -- 0x1200
    x"38",x"D0",x"F1",x"20",x"97",x"8A",x"C9",x"2C", -- 0x1208
    x"F0",x"03",x"4C",x"96",x"8B",x"4C",x"2F",x"91", -- 0x1210
    x"00",x"0B",x"DE",x"20",x"73",x"70",x"61",x"63", -- 0x1218
    x"65",x"00",x"E6",x"2A",x"D0",x"0A",x"E6",x"2B", -- 0x1220
    x"D0",x"06",x"E6",x"2C",x"D0",x"02",x"E6",x"2D", -- 0x1228
    x"60",x"A2",x"3F",x"20",x"0D",x"BE",x"A2",x"00", -- 0x1230
    x"A0",x"00",x"46",x"40",x"66",x"3F",x"90",x"0B", -- 0x1238
    x"18",x"98",x"65",x"2A",x"A8",x"8A",x"65",x"2B", -- 0x1240
    x"AA",x"B0",x"0F",x"06",x"2A",x"26",x"2B",x"A5", -- 0x1248
    x"3F",x"05",x"40",x"D0",x"E5",x"84",x"2A",x"86", -- 0x1250
    x"2B",x"60",x"4C",x"27",x"91",x"20",x"EB",x"92", -- 0x1258
    x"A5",x"2A",x"85",x"06",x"85",x"04",x"A5",x"2B", -- 0x1260
    x"85",x"07",x"85",x"05",x"4C",x"9B",x"8B",x"20", -- 0x1268
    x"EB",x"92",x"A5",x"2A",x"85",x"00",x"85",x"02", -- 0x1270
    x"A5",x"2B",x"85",x"01",x"85",x"03",x"20",x"2F", -- 0x1278
    x"BD",x"F0",x"07",x"20",x"EB",x"92",x"A5",x"2B", -- 0x1280
    x"85",x"18",x"4C",x"9B",x"8B",x"20",x"57",x"98", -- 0x1288
    x"20",x"20",x"BD",x"F0",x"F5",x"20",x"DF",x"97", -- 0x1290
    x"B0",x"0B",x"C9",x"EE",x"F0",x"19",x"C9",x"87", -- 0x1298
    x"F0",x"1E",x"20",x"21",x"88",x"20",x"57",x"98", -- 0x12A0
    x"A5",x"2A",x"85",x"21",x"A5",x"2B",x"85",x"22", -- 0x12A8
    x"A9",x"FF",x"85",x"20",x"4C",x"9B",x"8B",x"E6", -- 0x12B0
    x"0A",x"20",x"57",x"98",x"A9",x"FF",x"D0",x"EE", -- 0x12B8
    x"E6",x"0A",x"20",x"57",x"98",x"A9",x"00",x"F0", -- 0x12C0
    x"E9",x"20",x"EB",x"92",x"A2",x"2A",x"A0",x"00", -- 0x12C8
    x"84",x"2E",x"A9",x"02",x"20",x"F1",x"FF",x"4C", -- 0x12D0
    x"9B",x"8B",x"20",x"AE",x"8A",x"20",x"29",x"9B", -- 0x12D8
    x"4C",x"F0",x"92",x"20",x"EC",x"AD",x"F0",x"0F", -- 0x12E0
    x"30",x"0A",x"60",x"20",x"07",x"98",x"A5",x"27", -- 0x12E8
    x"F0",x"05",x"10",x"F6",x"4C",x"E4",x"A3",x"4C", -- 0x12F0
    x"0E",x"8C",x"20",x"EC",x"AD",x"F0",x"F8",x"30", -- 0x12F8
    x"E9",x"4C",x"BE",x"A2",x"A5",x"0B",x"85",x"19", -- 0x1300
    x"A5",x"0C",x"85",x"1A",x"A5",x"0A",x"85",x"1B", -- 0x1308
    x"A9",x"F2",x"20",x"97",x"B1",x"20",x"52",x"98", -- 0x1310
    x"4C",x"9B",x"8B",x"A0",x"03",x"A9",x"00",x"91", -- 0x1318
    x"2A",x"F0",x"1E",x"BA",x"E0",x"FC",x"B0",x"43", -- 0x1320
    x"20",x"82",x"95",x"F0",x"26",x"20",x"0D",x"B3", -- 0x1328
    x"A4",x"2C",x"30",x"E7",x"20",x"94",x"BD",x"A9", -- 0x1330
    x"00",x"20",x"D8",x"AE",x"85",x"27",x"20",x"B4", -- 0x1338
    x"B4",x"BA",x"FE",x"06",x"01",x"A4",x"1B",x"84", -- 0x1340
    x"0A",x"20",x"97",x"8A",x"C9",x"2C",x"F0",x"D3", -- 0x1348
    x"4C",x"96",x"8B",x"4C",x"98",x"8B",x"BA",x"E0", -- 0x1350
    x"FC",x"B0",x"0A",x"AD",x"FF",x"01",x"C9",x"F2", -- 0x1358
    x"D0",x"03",x"4C",x"57",x"98",x"00",x"0D",x"4E", -- 0x1360
    x"6F",x"20",x"F2",x"00",x"0C",x"4E",x"6F",x"74", -- 0x1368
    x"20",x"EA",x"00",x"19",x"42",x"61",x"64",x"20", -- 0x1370
    x"EB",x"00",x"20",x"21",x"88",x"A5",x"2A",x"48", -- 0x1378
    x"20",x"DA",x"92",x"20",x"52",x"98",x"A9",x"12", -- 0x1380
    x"20",x"EE",x"FF",x"4C",x"DA",x"93",x"A9",x"11", -- 0x1388
    x"48",x"20",x"21",x"88",x"20",x"57",x"98",x"4C", -- 0x1390
    x"DA",x"93",x"A9",x"16",x"48",x"20",x"21",x"88", -- 0x1398
    x"20",x"57",x"98",x"20",x"E7",x"BE",x"E0",x"FF", -- 0x13A0
    x"D0",x"2D",x"C0",x"FF",x"D0",x"29",x"A5",x"04", -- 0x13A8
    x"C5",x"06",x"D0",x"BE",x"A5",x"05",x"C5",x"07", -- 0x13B0
    x"D0",x"B8",x"A6",x"2A",x"A9",x"85",x"20",x"F4", -- 0x13B8
    x"FF",x"E4",x"02",x"98",x"E5",x"03",x"90",x"AA", -- 0x13C0
    x"E4",x"12",x"98",x"E5",x"13",x"90",x"A3",x"86", -- 0x13C8
    x"06",x"86",x"04",x"84",x"07",x"84",x"05",x"20", -- 0x13D0
    x"28",x"BC",x"68",x"20",x"EE",x"FF",x"20",x"56", -- 0x13D8
    x"94",x"4C",x"9B",x"8B",x"A9",x"04",x"D0",x"02", -- 0x13E0
    x"A9",x"05",x"48",x"20",x"1D",x"9B",x"4C",x"FD", -- 0x13E8
    x"93",x"20",x"21",x"88",x"A5",x"2A",x"48",x"20", -- 0x13F0
    x"AE",x"8A",x"20",x"29",x"9B",x"20",x"EE",x"92", -- 0x13F8
    x"20",x"94",x"BD",x"20",x"DA",x"92",x"20",x"52", -- 0x1400
    x"98",x"A9",x"19",x"20",x"EE",x"FF",x"68",x"20", -- 0x1408
    x"EE",x"FF",x"20",x"0B",x"BE",x"A5",x"37",x"20", -- 0x1410
    x"EE",x"FF",x"A5",x"38",x"20",x"EE",x"FF",x"20", -- 0x1418
    x"56",x"94",x"A5",x"2B",x"20",x"EE",x"FF",x"4C", -- 0x1420
    x"9B",x"8B",x"A5",x"2B",x"20",x"EE",x"FF",x"20", -- 0x1428
    x"97",x"8A",x"C9",x"3A",x"F0",x"1D",x"C9",x"0D", -- 0x1430
    x"F0",x"19",x"C9",x"8B",x"F0",x"15",x"C6",x"0A", -- 0x1438
    x"20",x"21",x"88",x"20",x"56",x"94",x"20",x"97", -- 0x1440
    x"8A",x"C9",x"2C",x"F0",x"E2",x"C9",x"3B",x"D0", -- 0x1448
    x"E1",x"F0",x"D7",x"4C",x"96",x"8B",x"A5",x"2A", -- 0x1450
    x"6C",x"0E",x"02",x"A0",x"01",x"B1",x"37",x"A0", -- 0x1458
    x"F6",x"C9",x"F2",x"F0",x"0A",x"A0",x"F8",x"D0", -- 0x1460
    x"06",x"A0",x"01",x"B1",x"37",x"0A",x"A8",x"B9", -- 0x1468
    x"00",x"04",x"85",x"3A",x"B9",x"01",x"04",x"85", -- 0x1470
    x"3B",x"A5",x"3B",x"F0",x"35",x"A0",x"00",x"B1", -- 0x1478
    x"3A",x"85",x"3C",x"C8",x"B1",x"3A",x"85",x"3D", -- 0x1480
    x"C8",x"B1",x"3A",x"D0",x"0D",x"88",x"C4",x"39", -- 0x1488
    x"D0",x"21",x"C8",x"B0",x"12",x"C8",x"B1",x"3A", -- 0x1490
    x"F0",x"19",x"D1",x"37",x"D0",x"15",x"C4",x"39", -- 0x1498
    x"D0",x"F3",x"C8",x"B1",x"3A",x"D0",x"0C",x"98", -- 0x14A0
    x"65",x"3A",x"85",x"2A",x"A5",x"3B",x"69",x"00", -- 0x14A8
    x"85",x"2B",x"60",x"A5",x"3D",x"F0",x"FB",x"A0", -- 0x14B0
    x"00",x"B1",x"3C",x"85",x"3A",x"C8",x"B1",x"3C", -- 0x14B8
    x"85",x"3B",x"C8",x"B1",x"3C",x"D0",x"0D",x"88", -- 0x14C0
    x"C4",x"39",x"D0",x"AD",x"C8",x"B0",x"12",x"C8", -- 0x14C8
    x"B1",x"3C",x"F0",x"A5",x"D1",x"37",x"D0",x"A1", -- 0x14D0
    x"C4",x"39",x"D0",x"F3",x"C8",x"B1",x"3C",x"D0", -- 0x14D8
    x"98",x"98",x"65",x"3C",x"85",x"2A",x"A5",x"3D", -- 0x14E0
    x"69",x"00",x"85",x"2B",x"60",x"A0",x"01",x"B1", -- 0x14E8
    x"37",x"AA",x"A9",x"F6",x"E0",x"F2",x"F0",x"09", -- 0x14F0
    x"A9",x"F8",x"D0",x"05",x"A0",x"01",x"B1",x"37", -- 0x14F8
    x"0A",x"85",x"3A",x"A9",x"04",x"85",x"3B",x"B1", -- 0x1500
    x"3A",x"F0",x"0B",x"AA",x"88",x"B1",x"3A",x"85", -- 0x1508
    x"3A",x"86",x"3B",x"C8",x"10",x"F1",x"A5",x"03", -- 0x1510
    x"91",x"3A",x"A5",x"02",x"88",x"91",x"3A",x"98", -- 0x1518
    x"C8",x"91",x"02",x"C4",x"39",x"F0",x"31",x"C8", -- 0x1520
    x"B1",x"37",x"91",x"02",x"C4",x"39",x"D0",x"F7", -- 0x1528
    x"60",x"A9",x"00",x"C8",x"91",x"02",x"CA",x"D0", -- 0x1530
    x"FA",x"38",x"98",x"65",x"02",x"90",x"02",x"E6", -- 0x1538
    x"03",x"A4",x"03",x"C4",x"05",x"90",x"0F",x"D0", -- 0x1540
    x"04",x"C5",x"04",x"90",x"09",x"A9",x"00",x"A0", -- 0x1548
    x"01",x"91",x"3A",x"4C",x"B7",x"8C",x"85",x"02", -- 0x1550
    x"60",x"A0",x"01",x"B1",x"37",x"C9",x"30",x"90", -- 0x1558
    x"18",x"C9",x"40",x"B0",x"0C",x"C9",x"3A",x"B0", -- 0x1560
    x"10",x"C0",x"01",x"F0",x"0C",x"E8",x"C8",x"D0", -- 0x1568
    x"EA",x"C9",x"5F",x"B0",x"05",x"C9",x"5B",x"90", -- 0x1570
    x"F4",x"60",x"C9",x"7B",x"90",x"EF",x"60",x"20", -- 0x1578
    x"31",x"95",x"20",x"C9",x"95",x"D0",x"1D",x"B0", -- 0x1580
    x"1B",x"20",x"FC",x"94",x"A2",x"05",x"E4",x"2C", -- 0x1588
    x"D0",x"ED",x"E8",x"D0",x"EA",x"C9",x"21",x"F0", -- 0x1590
    x"0C",x"C9",x"24",x"F0",x"13",x"49",x"3F",x"F0", -- 0x1598
    x"06",x"A9",x"00",x"38",x"60",x"A9",x"04",x"48", -- 0x15A0
    x"E6",x"1B",x"20",x"E3",x"92",x"4C",x"9F",x"96", -- 0x15A8
    x"E6",x"1B",x"20",x"E3",x"92",x"A5",x"2B",x"F0", -- 0x15B0
    x"06",x"A9",x"80",x"85",x"2C",x"38",x"60",x"00", -- 0x15B8
    x"08",x"24",x"20",x"72",x"61",x"6E",x"67",x"65", -- 0x15C0
    x"00",x"A5",x"0B",x"85",x"19",x"A5",x"0C",x"85", -- 0x15C8
    x"1A",x"A4",x"0A",x"88",x"C8",x"84",x"1B",x"B1", -- 0x15D0
    x"19",x"C9",x"20",x"F0",x"F7",x"C9",x"40",x"90", -- 0x15D8
    x"B4",x"C9",x"5B",x"B0",x"1A",x"0A",x"0A",x"85", -- 0x15E0
    x"2A",x"A9",x"04",x"85",x"2B",x"C8",x"B1",x"19", -- 0x15E8
    x"C8",x"C9",x"25",x"D0",x"0A",x"A2",x"04",x"86", -- 0x15F0
    x"2C",x"B1",x"19",x"C9",x"28",x"D0",x"66",x"A2", -- 0x15F8
    x"05",x"86",x"2C",x"A5",x"1B",x"18",x"65",x"19", -- 0x1600
    x"A6",x"1A",x"90",x"02",x"E8",x"18",x"E9",x"00", -- 0x1608
    x"85",x"37",x"B0",x"01",x"CA",x"86",x"38",x"A6", -- 0x1610
    x"1B",x"A0",x"01",x"B1",x"37",x"C9",x"41",x"B0", -- 0x1618
    x"0C",x"C9",x"30",x"90",x"1C",x"C9",x"3A",x"B0", -- 0x1620
    x"18",x"E8",x"C8",x"D0",x"EE",x"C9",x"5B",x"B0", -- 0x1628
    x"04",x"E8",x"C8",x"D0",x"E6",x"C9",x"5F",x"90", -- 0x1630
    x"08",x"C9",x"7B",x"B0",x"04",x"E8",x"C8",x"D0", -- 0x1638
    x"DA",x"88",x"F0",x"2F",x"C9",x"24",x"F0",x"67", -- 0x1640
    x"C9",x"25",x"D0",x"08",x"C6",x"2C",x"C8",x"E8", -- 0x1648
    x"C8",x"B1",x"37",x"88",x"84",x"39",x"C9",x"28", -- 0x1650
    x"F0",x"4C",x"20",x"69",x"94",x"F0",x"18",x"86", -- 0x1658
    x"1B",x"A4",x"1B",x"B1",x"19",x"C9",x"21",x"F0", -- 0x1660
    x"16",x"C9",x"3F",x"F0",x"0E",x"18",x"84",x"1B", -- 0x1668
    x"A9",x"FF",x"60",x"A9",x"00",x"38",x"60",x"A9", -- 0x1670
    x"00",x"18",x"60",x"A9",x"00",x"F0",x"02",x"A9", -- 0x1678
    x"04",x"48",x"C8",x"84",x"1B",x"20",x"2C",x"B3", -- 0x1680
    x"20",x"F0",x"92",x"A5",x"2B",x"48",x"A5",x"2A", -- 0x1688
    x"48",x"20",x"E3",x"92",x"18",x"68",x"65",x"2A", -- 0x1690
    x"85",x"2A",x"68",x"65",x"2B",x"85",x"2B",x"68", -- 0x1698
    x"85",x"2C",x"18",x"A9",x"FF",x"60",x"E8",x"E6", -- 0x16A0
    x"39",x"20",x"DF",x"96",x"4C",x"61",x"96",x"E8", -- 0x16A8
    x"C8",x"84",x"39",x"C8",x"C6",x"2C",x"B1",x"37", -- 0x16B0
    x"C9",x"28",x"F0",x"0D",x"20",x"69",x"94",x"F0", -- 0x16B8
    x"B6",x"86",x"1B",x"A9",x"81",x"85",x"2C",x"38", -- 0x16C0
    x"60",x"E8",x"84",x"39",x"C6",x"2C",x"20",x"DF", -- 0x16C8
    x"96",x"A9",x"81",x"85",x"2C",x"38",x"60",x"00", -- 0x16D0
    x"0E",x"41",x"72",x"72",x"61",x"79",x"00",x"20", -- 0x16D8
    x"69",x"94",x"F0",x"F3",x"86",x"1B",x"A5",x"2C", -- 0x16E0
    x"48",x"A5",x"2A",x"48",x"A5",x"2B",x"48",x"A0", -- 0x16E8
    x"00",x"B1",x"2A",x"C9",x"04",x"90",x"75",x"98", -- 0x16F0
    x"20",x"D8",x"AE",x"A9",x"01",x"85",x"2D",x"20", -- 0x16F8
    x"94",x"BD",x"20",x"DD",x"92",x"E6",x"1B",x"E0", -- 0x1700
    x"2C",x"D0",x"CC",x"A2",x"39",x"20",x"0D",x"BE", -- 0x1708
    x"A4",x"3C",x"68",x"85",x"38",x"68",x"85",x"37", -- 0x1710
    x"48",x"A5",x"38",x"48",x"20",x"BA",x"97",x"84", -- 0x1718
    x"2D",x"B1",x"37",x"85",x"3F",x"C8",x"B1",x"37", -- 0x1720
    x"85",x"40",x"A5",x"2A",x"65",x"39",x"85",x"2A", -- 0x1728
    x"A5",x"2B",x"65",x"3A",x"85",x"2B",x"20",x"36", -- 0x1730
    x"92",x"A0",x"00",x"38",x"B1",x"37",x"E5",x"2D", -- 0x1738
    x"C9",x"03",x"B0",x"BB",x"20",x"94",x"BD",x"20", -- 0x1740
    x"56",x"AE",x"20",x"F0",x"92",x"68",x"85",x"38", -- 0x1748
    x"68",x"85",x"37",x"A2",x"39",x"20",x"0D",x"BE", -- 0x1750
    x"A4",x"3C",x"20",x"BA",x"97",x"18",x"A5",x"39", -- 0x1758
    x"65",x"2A",x"85",x"2A",x"A5",x"3A",x"65",x"2B", -- 0x1760
    x"85",x"2B",x"90",x"11",x"20",x"56",x"AE",x"20", -- 0x1768
    x"F0",x"92",x"68",x"85",x"38",x"68",x"85",x"37", -- 0x1770
    x"A0",x"01",x"20",x"BA",x"97",x"68",x"85",x"2C", -- 0x1778
    x"C9",x"05",x"D0",x"17",x"A6",x"2B",x"A5",x"2A", -- 0x1780
    x"06",x"2A",x"26",x"2B",x"06",x"2A",x"26",x"2B", -- 0x1788
    x"65",x"2A",x"85",x"2A",x"8A",x"65",x"2B",x"85", -- 0x1790
    x"2B",x"90",x"08",x"06",x"2A",x"26",x"2B",x"06", -- 0x1798
    x"2A",x"26",x"2B",x"98",x"65",x"2A",x"85",x"2A", -- 0x17A0
    x"90",x"03",x"E6",x"2B",x"18",x"A5",x"37",x"65", -- 0x17A8
    x"2A",x"85",x"2A",x"A5",x"38",x"65",x"2B",x"85", -- 0x17B0
    x"2B",x"60",x"A5",x"2B",x"29",x"C0",x"05",x"2C", -- 0x17B8
    x"05",x"2D",x"D0",x"0D",x"A5",x"2A",x"D1",x"37", -- 0x17C0
    x"C8",x"A5",x"2B",x"F1",x"37",x"B0",x"02",x"C8", -- 0x17C8
    x"60",x"00",x"0F",x"53",x"75",x"62",x"73",x"63", -- 0x17D0
    x"72",x"69",x"70",x"74",x"00",x"E6",x"0A",x"A4", -- 0x17D8
    x"0A",x"B1",x"0B",x"C9",x"20",x"F0",x"F6",x"C9", -- 0x17E0
    x"8D",x"D0",x"1A",x"C8",x"B1",x"0B",x"0A",x"0A", -- 0x17E8
    x"AA",x"29",x"C0",x"C8",x"51",x"0B",x"85",x"2A", -- 0x17F0
    x"8A",x"0A",x"0A",x"C8",x"51",x"0B",x"85",x"2B", -- 0x17F8
    x"C8",x"84",x"0A",x"38",x"60",x"18",x"60",x"A5", -- 0x1800
    x"0B",x"85",x"19",x"A5",x"0C",x"85",x"1A",x"A5", -- 0x1808
    x"0A",x"85",x"1B",x"A4",x"1B",x"E6",x"1B",x"B1", -- 0x1810
    x"19",x"C9",x"20",x"F0",x"F6",x"C9",x"3D",x"F0", -- 0x1818
    x"28",x"00",x"04",x"4D",x"69",x"73",x"74",x"61", -- 0x1820
    x"6B",x"65",x"00",x"10",x"53",x"79",x"6E",x"74", -- 0x1828
    x"61",x"78",x"20",x"65",x"72",x"72",x"6F",x"72", -- 0x1830
    x"00",x"11",x"45",x"73",x"63",x"61",x"70",x"65", -- 0x1838
    x"00",x"20",x"8C",x"8A",x"C9",x"3D",x"D0",x"D9", -- 0x1840
    x"60",x"20",x"29",x"9B",x"8A",x"A4",x"1B",x"4C", -- 0x1848
    x"61",x"98",x"A4",x"1B",x"4C",x"59",x"98",x"A4", -- 0x1850
    x"0A",x"88",x"C8",x"B1",x"0B",x"C9",x"20",x"F0", -- 0x1858
    x"F9",x"C9",x"3A",x"F0",x"08",x"C9",x"0D",x"F0", -- 0x1860
    x"04",x"C9",x"8B",x"D0",x"BD",x"18",x"98",x"65", -- 0x1868
    x"0B",x"85",x"0B",x"90",x"02",x"E6",x"0C",x"A0", -- 0x1870
    x"01",x"84",x"0A",x"24",x"FF",x"30",x"B9",x"60", -- 0x1878
    x"20",x"57",x"98",x"88",x"B1",x"0B",x"C9",x"3A", -- 0x1880
    x"F0",x"F5",x"A5",x"0C",x"C9",x"07",x"F0",x"2C", -- 0x1888
    x"C8",x"B1",x"0B",x"30",x"27",x"A5",x"20",x"F0", -- 0x1890
    x"13",x"98",x"48",x"C8",x"B1",x"0B",x"48",x"88", -- 0x1898
    x"B1",x"0B",x"A8",x"68",x"20",x"EA",x"AE",x"20", -- 0x18A0
    x"05",x"99",x"68",x"A8",x"C8",x"38",x"98",x"65", -- 0x18A8
    x"0B",x"85",x"0B",x"90",x"02",x"E6",x"0C",x"A0", -- 0x18B0
    x"01",x"84",x"0A",x"60",x"4C",x"F6",x"8A",x"4C", -- 0x18B8
    x"0E",x"8C",x"20",x"1D",x"9B",x"F0",x"F8",x"10", -- 0x18C0
    x"03",x"20",x"E4",x"A3",x"A4",x"1B",x"84",x"0A", -- 0x18C8
    x"A5",x"2A",x"05",x"2B",x"05",x"2C",x"05",x"2D", -- 0x18D0
    x"F0",x"17",x"E0",x"8C",x"F0",x"03",x"4C",x"A3", -- 0x18D8
    x"8B",x"E6",x"0A",x"20",x"DF",x"97",x"90",x"F6", -- 0x18E0
    x"20",x"AF",x"B9",x"20",x"77",x"98",x"4C",x"D2", -- 0x18E8
    x"B8",x"A4",x"0A",x"B1",x"0B",x"C9",x"0D",x"F0", -- 0x18F0
    x"09",x"C8",x"C9",x"8B",x"D0",x"F5",x"84",x"0A", -- 0x18F8
    x"F0",x"E1",x"4C",x"87",x"8B",x"A5",x"2A",x"C5", -- 0x1900
    x"21",x"A5",x"2B",x"E5",x"22",x"B0",x"AC",x"A9", -- 0x1908
    x"5B",x"20",x"58",x"B5",x"20",x"1F",x"99",x"A9", -- 0x1910
    x"5D",x"20",x"58",x"B5",x"4C",x"65",x"B5",x"A9", -- 0x1918
    x"00",x"F0",x"02",x"A9",x"05",x"85",x"14",x"A2", -- 0x1920
    x"04",x"A9",x"00",x"95",x"3F",x"38",x"A5",x"2A", -- 0x1928
    x"FD",x"6B",x"99",x"A8",x"A5",x"2B",x"FD",x"B9", -- 0x1930
    x"99",x"90",x"08",x"85",x"2B",x"84",x"2A",x"F6", -- 0x1938
    x"3F",x"D0",x"EB",x"CA",x"10",x"E3",x"A2",x"05", -- 0x1940
    x"CA",x"F0",x"04",x"B5",x"3F",x"F0",x"F9",x"86", -- 0x1948
    x"37",x"A5",x"14",x"F0",x"0B",x"E5",x"37",x"F0", -- 0x1950
    x"07",x"A8",x"20",x"65",x"B5",x"88",x"D0",x"FA", -- 0x1958
    x"B5",x"3F",x"09",x"30",x"20",x"58",x"B5",x"CA", -- 0x1960
    x"10",x"F6",x"60",x"01",x"0A",x"64",x"E8",x"10", -- 0x1968
    x"A0",x"00",x"84",x"3D",x"A5",x"18",x"85",x"3E", -- 0x1970
    x"A0",x"01",x"B1",x"3D",x"C5",x"2B",x"B0",x"0E", -- 0x1978
    x"A0",x"03",x"B1",x"3D",x"65",x"3D",x"85",x"3D", -- 0x1980
    x"90",x"EE",x"E6",x"3E",x"B0",x"EA",x"D0",x"14", -- 0x1988
    x"A0",x"02",x"B1",x"3D",x"C5",x"2A",x"90",x"E8", -- 0x1990
    x"D0",x"0A",x"98",x"65",x"3D",x"85",x"3D",x"90", -- 0x1998
    x"03",x"E6",x"3E",x"18",x"A0",x"02",x"60",x"00", -- 0x19A0
    x"12",x"44",x"69",x"76",x"69",x"73",x"69",x"6F", -- 0x19A8
    x"6E",x"20",x"62",x"79",x"20",x"7A",x"65",x"72", -- 0x19B0
    x"6F",x"00",x"00",x"00",x"03",x"27",x"A8",x"20", -- 0x19B8
    x"F0",x"92",x"A5",x"2D",x"48",x"20",x"71",x"AD", -- 0x19C0
    x"20",x"1D",x"9E",x"86",x"27",x"A8",x"20",x"F0", -- 0x19C8
    x"92",x"68",x"85",x"38",x"45",x"2D",x"85",x"37", -- 0x19D0
    x"20",x"71",x"AD",x"A2",x"39",x"20",x"0D",x"BE", -- 0x19D8
    x"84",x"3D",x"84",x"3E",x"84",x"3F",x"84",x"40", -- 0x19E0
    x"A5",x"2D",x"05",x"2A",x"05",x"2B",x"05",x"2C", -- 0x19E8
    x"F0",x"B5",x"A0",x"20",x"88",x"F0",x"41",x"06", -- 0x19F0
    x"39",x"26",x"3A",x"26",x"3B",x"26",x"3C",x"10", -- 0x19F8
    x"F3",x"26",x"39",x"26",x"3A",x"26",x"3B",x"26", -- 0x1A00
    x"3C",x"26",x"3D",x"26",x"3E",x"26",x"3F",x"26", -- 0x1A08
    x"40",x"38",x"A5",x"3D",x"E5",x"2A",x"48",x"A5", -- 0x1A10
    x"3E",x"E5",x"2B",x"48",x"A5",x"3F",x"E5",x"2C", -- 0x1A18
    x"AA",x"A5",x"40",x"E5",x"2D",x"90",x"0C",x"85", -- 0x1A20
    x"40",x"86",x"3F",x"68",x"85",x"3E",x"68",x"85", -- 0x1A28
    x"3D",x"B0",x"02",x"68",x"68",x"88",x"D0",x"C9", -- 0x1A30
    x"60",x"86",x"27",x"20",x"EA",x"BD",x"20",x"51", -- 0x1A38
    x"BD",x"20",x"BE",x"A2",x"20",x"1E",x"A2",x"20", -- 0x1A40
    x"7E",x"BD",x"20",x"B5",x"A3",x"4C",x"62",x"9A", -- 0x1A48
    x"20",x"51",x"BD",x"20",x"42",x"9C",x"86",x"27", -- 0x1A50
    x"A8",x"20",x"FD",x"92",x"20",x"7E",x"BD",x"20", -- 0x1A58
    x"4E",x"A3",x"A6",x"27",x"A0",x"00",x"A5",x"3B", -- 0x1A60
    x"29",x"80",x"85",x"3B",x"A5",x"2E",x"29",x"80", -- 0x1A68
    x"C5",x"3B",x"D0",x"1E",x"A5",x"3D",x"C5",x"30", -- 0x1A70
    x"D0",x"19",x"A5",x"3E",x"C5",x"31",x"D0",x"13", -- 0x1A78
    x"A5",x"3F",x"C5",x"32",x"D0",x"0D",x"A5",x"40", -- 0x1A80
    x"C5",x"33",x"D0",x"07",x"A5",x"41",x"C5",x"34", -- 0x1A88
    x"D0",x"01",x"60",x"6A",x"45",x"3B",x"2A",x"A9", -- 0x1A90
    x"01",x"60",x"4C",x"0E",x"8C",x"8A",x"F0",x"47", -- 0x1A98
    x"30",x"AE",x"20",x"94",x"BD",x"20",x"42",x"9C", -- 0x1AA0
    x"A8",x"F0",x"EF",x"30",x"8C",x"A5",x"2D",x"49", -- 0x1AA8
    x"80",x"85",x"2D",x"38",x"A0",x"00",x"B1",x"04", -- 0x1AB0
    x"E5",x"2A",x"85",x"2A",x"C8",x"B1",x"04",x"E5", -- 0x1AB8
    x"2B",x"85",x"2B",x"C8",x"B1",x"04",x"E5",x"2C", -- 0x1AC0
    x"85",x"2C",x"C8",x"B1",x"04",x"A0",x"00",x"49", -- 0x1AC8
    x"80",x"E5",x"2D",x"05",x"2A",x"05",x"2B",x"05", -- 0x1AD0
    x"2C",x"08",x"18",x"A9",x"04",x"65",x"04",x"85", -- 0x1AD8
    x"04",x"90",x"02",x"E6",x"05",x"28",x"60",x"20", -- 0x1AE0
    x"B2",x"BD",x"20",x"42",x"9C",x"A8",x"D0",x"AA", -- 0x1AE8
    x"86",x"37",x"A6",x"36",x"A0",x"00",x"B1",x"04", -- 0x1AF0
    x"85",x"39",x"C5",x"36",x"B0",x"01",x"AA",x"86", -- 0x1AF8
    x"3A",x"A0",x"00",x"C4",x"3A",x"F0",x"0A",x"C8", -- 0x1B00
    x"B1",x"04",x"D9",x"FF",x"05",x"F0",x"F4",x"D0", -- 0x1B08
    x"04",x"A5",x"39",x"C5",x"36",x"08",x"20",x"DC", -- 0x1B10
    x"BD",x"A6",x"37",x"28",x"60",x"A5",x"0B",x"85", -- 0x1B18
    x"19",x"A5",x"0C",x"85",x"1A",x"A5",x"0A",x"85", -- 0x1B20
    x"1B",x"20",x"72",x"9B",x"E0",x"84",x"F0",x"0A", -- 0x1B28
    x"E0",x"82",x"F0",x"21",x"C6",x"1B",x"A8",x"85", -- 0x1B30
    x"27",x"60",x"20",x"6B",x"9B",x"A8",x"20",x"F0", -- 0x1B38
    x"92",x"A0",x"03",x"B1",x"04",x"19",x"2A",x"00", -- 0x1B40
    x"99",x"2A",x"00",x"88",x"10",x"F5",x"20",x"FF", -- 0x1B48
    x"BD",x"A9",x"40",x"D0",x"D7",x"20",x"6B",x"9B", -- 0x1B50
    x"A8",x"20",x"F0",x"92",x"A0",x"03",x"B1",x"04", -- 0x1B58
    x"59",x"2A",x"00",x"99",x"2A",x"00",x"88",x"10", -- 0x1B60
    x"F5",x"30",x"E3",x"A8",x"20",x"F0",x"92",x"20", -- 0x1B68
    x"94",x"BD",x"20",x"9C",x"9B",x"E0",x"80",x"F0", -- 0x1B70
    x"01",x"60",x"A8",x"20",x"F0",x"92",x"20",x"94", -- 0x1B78
    x"BD",x"20",x"9C",x"9B",x"A8",x"20",x"F0",x"92", -- 0x1B80
    x"A0",x"03",x"B1",x"04",x"39",x"2A",x"00",x"99", -- 0x1B88
    x"2A",x"00",x"88",x"10",x"F5",x"20",x"FF",x"BD", -- 0x1B90
    x"A9",x"40",x"D0",x"D9",x"20",x"42",x"9C",x"E0", -- 0x1B98
    x"3F",x"B0",x"04",x"E0",x"3C",x"B0",x"01",x"60", -- 0x1BA0
    x"F0",x"16",x"E0",x"3E",x"F0",x"3A",x"AA",x"20", -- 0x1BA8
    x"9E",x"9A",x"D0",x"01",x"88",x"84",x"2A",x"84", -- 0x1BB0
    x"2B",x"84",x"2C",x"84",x"2D",x"A9",x"40",x"60", -- 0x1BB8
    x"AA",x"A4",x"1B",x"B1",x"19",x"C9",x"3D",x"F0", -- 0x1BC0
    x"0B",x"C9",x"3E",x"F0",x"12",x"20",x"9D",x"9A", -- 0x1BC8
    x"90",x"E2",x"B0",x"E1",x"E6",x"1B",x"20",x"9D", -- 0x1BD0
    x"9A",x"F0",x"D9",x"90",x"D7",x"B0",x"D6",x"E6", -- 0x1BD8
    x"1B",x"20",x"9D",x"9A",x"D0",x"CE",x"F0",x"CD", -- 0x1BE0
    x"AA",x"A4",x"1B",x"B1",x"19",x"C9",x"3D",x"F0", -- 0x1BE8
    x"09",x"20",x"9D",x"9A",x"F0",x"BF",x"B0",x"BC", -- 0x1BF0
    x"90",x"BB",x"E6",x"1B",x"20",x"9D",x"9A",x"B0", -- 0x1BF8
    x"B3",x"90",x"B2",x"00",x"13",x"53",x"74",x"72", -- 0x1C00
    x"69",x"6E",x"67",x"20",x"74",x"6F",x"6F",x"20", -- 0x1C08
    x"6C",x"6F",x"6E",x"67",x"00",x"20",x"B2",x"BD", -- 0x1C10
    x"20",x"20",x"9E",x"A8",x"D0",x"6A",x"18",x"86", -- 0x1C18
    x"37",x"A0",x"00",x"B1",x"04",x"65",x"36",x"B0", -- 0x1C20
    x"DA",x"AA",x"48",x"A4",x"36",x"B9",x"FF",x"05", -- 0x1C28
    x"9D",x"FF",x"05",x"CA",x"88",x"D0",x"F6",x"20", -- 0x1C30
    x"CB",x"BD",x"68",x"85",x"36",x"A6",x"37",x"98", -- 0x1C38
    x"F0",x"03",x"20",x"D1",x"9D",x"E0",x"2B",x"F0", -- 0x1C40
    x"05",x"E0",x"2D",x"F0",x"68",x"60",x"A8",x"F0", -- 0x1C48
    x"C4",x"30",x"38",x"20",x"CE",x"9D",x"A8",x"F0", -- 0x1C50
    x"2F",x"30",x"4C",x"A0",x"00",x"18",x"B1",x"04", -- 0x1C58
    x"65",x"2A",x"85",x"2A",x"C8",x"B1",x"04",x"65", -- 0x1C60
    x"2B",x"85",x"2B",x"C8",x"B1",x"04",x"65",x"2C", -- 0x1C68
    x"85",x"2C",x"C8",x"B1",x"04",x"65",x"2D",x"85", -- 0x1C70
    x"2D",x"18",x"A5",x"04",x"69",x"04",x"85",x"04", -- 0x1C78
    x"A9",x"40",x"90",x"C1",x"E6",x"05",x"B0",x"BD", -- 0x1C80
    x"4C",x"0E",x"8C",x"20",x"51",x"BD",x"20",x"D1", -- 0x1C88
    x"9D",x"A8",x"F0",x"F4",x"86",x"27",x"30",x"03", -- 0x1C90
    x"20",x"BE",x"A2",x"20",x"7E",x"BD",x"20",x"00", -- 0x1C98
    x"A5",x"A6",x"27",x"A9",x"FF",x"D0",x"9E",x"86", -- 0x1CA0
    x"27",x"20",x"EA",x"BD",x"20",x"51",x"BD",x"20", -- 0x1CA8
    x"BE",x"A2",x"4C",x"9B",x"9C",x"A8",x"F0",x"D0", -- 0x1CB0
    x"30",x"27",x"20",x"CE",x"9D",x"A8",x"F0",x"C8", -- 0x1CB8
    x"30",x"38",x"38",x"A0",x"00",x"B1",x"04",x"E5", -- 0x1CC0
    x"2A",x"85",x"2A",x"C8",x"B1",x"04",x"E5",x"2B", -- 0x1CC8
    x"85",x"2B",x"C8",x"B1",x"04",x"E5",x"2C",x"85", -- 0x1CD0
    x"2C",x"C8",x"B1",x"04",x"E5",x"2D",x"4C",x"77", -- 0x1CD8
    x"9C",x"20",x"51",x"BD",x"20",x"D1",x"9D",x"A8", -- 0x1CE0
    x"F0",x"9E",x"86",x"27",x"30",x"03",x"20",x"BE", -- 0x1CE8
    x"A2",x"20",x"7E",x"BD",x"20",x"FD",x"A4",x"4C", -- 0x1CF0
    x"A1",x"9C",x"86",x"27",x"20",x"EA",x"BD",x"20", -- 0x1CF8
    x"51",x"BD",x"20",x"BE",x"A2",x"20",x"7E",x"BD", -- 0x1D00
    x"20",x"D0",x"A4",x"4C",x"A1",x"9C",x"20",x"BE", -- 0x1D08
    x"A2",x"20",x"EA",x"BD",x"20",x"51",x"BD",x"20", -- 0x1D10
    x"BE",x"A2",x"4C",x"2C",x"9D",x"20",x"BE",x"A2", -- 0x1D18
    x"20",x"51",x"BD",x"20",x"20",x"9E",x"86",x"27", -- 0x1D20
    x"A8",x"20",x"FD",x"92",x"20",x"7E",x"BD",x"20", -- 0x1D28
    x"56",x"A6",x"A9",x"FF",x"A6",x"27",x"4C",x"D4", -- 0x1D30
    x"9D",x"4C",x"0E",x"8C",x"A8",x"F0",x"FA",x"30", -- 0x1D38
    x"DF",x"A5",x"2D",x"C5",x"2C",x"D0",x"D6",x"A8", -- 0x1D40
    x"F0",x"04",x"C9",x"FF",x"D0",x"CF",x"45",x"2B", -- 0x1D48
    x"30",x"CB",x"20",x"1D",x"9E",x"86",x"27",x"A8", -- 0x1D50
    x"F0",x"DF",x"30",x"B5",x"A5",x"2D",x"C5",x"2C", -- 0x1D58
    x"D0",x"AC",x"A8",x"F0",x"04",x"C9",x"FF",x"D0", -- 0x1D60
    x"A5",x"45",x"2B",x"30",x"A1",x"A5",x"2D",x"48", -- 0x1D68
    x"20",x"71",x"AD",x"A2",x"39",x"20",x"44",x"BE", -- 0x1D70
    x"20",x"EA",x"BD",x"68",x"45",x"2D",x"85",x"37", -- 0x1D78
    x"20",x"71",x"AD",x"A0",x"00",x"A2",x"00",x"84", -- 0x1D80
    x"3F",x"84",x"40",x"46",x"3A",x"66",x"39",x"90", -- 0x1D88
    x"15",x"18",x"98",x"65",x"2A",x"A8",x"8A",x"65", -- 0x1D90
    x"2B",x"AA",x"A5",x"3F",x"65",x"2C",x"85",x"3F", -- 0x1D98
    x"A5",x"40",x"65",x"2D",x"85",x"40",x"06",x"2A", -- 0x1DA0
    x"26",x"2B",x"26",x"2C",x"26",x"2D",x"A5",x"39", -- 0x1DA8
    x"05",x"3A",x"D0",x"D7",x"84",x"3D",x"86",x"3E", -- 0x1DB0
    x"A5",x"37",x"08",x"A2",x"3D",x"20",x"56",x"AF", -- 0x1DB8
    x"28",x"10",x"03",x"20",x"93",x"AD",x"A6",x"27", -- 0x1DC0
    x"4C",x"D4",x"9D",x"4C",x"3C",x"9D",x"20",x"94", -- 0x1DC8
    x"BD",x"20",x"20",x"9E",x"E0",x"2A",x"F0",x"F3", -- 0x1DD0
    x"E0",x"2F",x"F0",x"09",x"E0",x"83",x"F0",x"21", -- 0x1DD8
    x"E0",x"81",x"F0",x"26",x"60",x"A8",x"20",x"FD", -- 0x1DE0
    x"92",x"20",x"51",x"BD",x"20",x"20",x"9E",x"86", -- 0x1DE8
    x"27",x"A8",x"20",x"FD",x"92",x"20",x"7E",x"BD", -- 0x1DF0
    x"20",x"AD",x"A6",x"A6",x"27",x"A9",x"FF",x"D0", -- 0x1DF8
    x"D3",x"20",x"BE",x"99",x"A5",x"38",x"08",x"4C", -- 0x1E00
    x"BB",x"9D",x"20",x"BE",x"99",x"26",x"39",x"26", -- 0x1E08
    x"3A",x"26",x"3B",x"26",x"3C",x"24",x"37",x"08", -- 0x1E10
    x"A2",x"39",x"4C",x"BD",x"9D",x"20",x"94",x"BD", -- 0x1E18
    x"20",x"EC",x"AD",x"48",x"A4",x"1B",x"E6",x"1B", -- 0x1E20
    x"B1",x"19",x"C9",x"20",x"F0",x"F6",x"AA",x"68", -- 0x1E28
    x"E0",x"5E",x"F0",x"01",x"60",x"A8",x"20",x"FD", -- 0x1E30
    x"92",x"20",x"51",x"BD",x"20",x"FA",x"92",x"A5", -- 0x1E38
    x"30",x"C9",x"87",x"B0",x"43",x"20",x"86",x"A4", -- 0x1E40
    x"D0",x"0F",x"20",x"7E",x"BD",x"20",x"B5",x"A3", -- 0x1E48
    x"A5",x"4A",x"20",x"12",x"AB",x"A9",x"FF",x"D0", -- 0x1E50
    x"CA",x"20",x"81",x"A3",x"A5",x"04",x"85",x"4B", -- 0x1E58
    x"A5",x"05",x"85",x"4C",x"20",x"B5",x"A3",x"A5", -- 0x1E60
    x"4A",x"20",x"12",x"AB",x"20",x"7D",x"A3",x"20", -- 0x1E68
    x"7E",x"BD",x"20",x"B5",x"A3",x"20",x"01",x"A8", -- 0x1E70
    x"20",x"D1",x"AA",x"20",x"94",x"AA",x"20",x"ED", -- 0x1E78
    x"A7",x"20",x"56",x"A6",x"A9",x"FF",x"D0",x"9B", -- 0x1E80
    x"20",x"81",x"A3",x"20",x"99",x"A6",x"D0",x"DC", -- 0x1E88
    x"98",x"10",x"03",x"20",x"E4",x"A3",x"A2",x"00", -- 0x1E90
    x"A0",x"00",x"B9",x"2A",x"00",x"48",x"29",x"0F", -- 0x1E98
    x"95",x"3F",x"68",x"4A",x"4A",x"4A",x"4A",x"E8", -- 0x1EA0
    x"95",x"3F",x"E8",x"C8",x"C0",x"04",x"D0",x"EA", -- 0x1EA8
    x"CA",x"F0",x"04",x"B5",x"3F",x"F0",x"F9",x"B5", -- 0x1EB0
    x"3F",x"C9",x"0A",x"90",x"02",x"69",x"06",x"69", -- 0x1EB8
    x"30",x"20",x"66",x"A0",x"CA",x"10",x"F0",x"60", -- 0x1EC0
    x"10",x"07",x"A9",x"2D",x"85",x"2E",x"20",x"66", -- 0x1EC8
    x"A0",x"A5",x"30",x"C9",x"81",x"B0",x"4E",x"20", -- 0x1ED0
    x"F4",x"A1",x"C6",x"49",x"4C",x"D1",x"9E",x"AE", -- 0x1ED8
    x"02",x"04",x"E0",x"03",x"90",x"02",x"A2",x"00", -- 0x1EE0
    x"86",x"37",x"AD",x"01",x"04",x"F0",x"06",x"C9", -- 0x1EE8
    x"0A",x"B0",x"06",x"90",x"06",x"E0",x"02",x"F0", -- 0x1EF0
    x"02",x"A9",x"0A",x"85",x"38",x"85",x"4E",x"A9", -- 0x1EF8
    x"00",x"85",x"36",x"85",x"49",x"24",x"15",x"30", -- 0x1F00
    x"87",x"98",x"30",x"03",x"20",x"BE",x"A2",x"20", -- 0x1F08
    x"DA",x"A1",x"D0",x"B4",x"A5",x"37",x"D0",x"05", -- 0x1F10
    x"A9",x"30",x"4C",x"66",x"A0",x"4C",x"9C",x"9F", -- 0x1F18
    x"20",x"99",x"A6",x"D0",x"0F",x"C9",x"84",x"90", -- 0x1F20
    x"10",x"D0",x"06",x"A5",x"31",x"C9",x"A0",x"90", -- 0x1F28
    x"08",x"20",x"4D",x"A2",x"E6",x"49",x"4C",x"D1", -- 0x1F30
    x"9E",x"A5",x"35",x"85",x"27",x"20",x"85",x"A3", -- 0x1F38
    x"A5",x"4E",x"85",x"38",x"A6",x"37",x"E0",x"02", -- 0x1F40
    x"D0",x"12",x"65",x"49",x"30",x"52",x"85",x"38", -- 0x1F48
    x"C9",x"0B",x"90",x"08",x"A9",x"0A",x"85",x"38", -- 0x1F50
    x"A9",x"00",x"85",x"37",x"20",x"86",x"A6",x"A9", -- 0x1F58
    x"A0",x"85",x"31",x"A9",x"83",x"85",x"30",x"A6", -- 0x1F60
    x"38",x"F0",x"06",x"20",x"4D",x"A2",x"CA",x"D0", -- 0x1F68
    x"FA",x"20",x"F5",x"A7",x"20",x"4E",x"A3",x"A5", -- 0x1F70
    x"27",x"85",x"42",x"20",x"0B",x"A5",x"A5",x"30", -- 0x1F78
    x"C9",x"84",x"B0",x"0E",x"66",x"31",x"66",x"32", -- 0x1F80
    x"66",x"33",x"66",x"34",x"66",x"35",x"E6",x"30", -- 0x1F88
    x"D0",x"EC",x"A5",x"31",x"C9",x"A0",x"B0",x"88", -- 0x1F90
    x"A5",x"38",x"D0",x"11",x"C9",x"01",x"F0",x"46", -- 0x1F98
    x"20",x"86",x"A6",x"A9",x"00",x"85",x"49",x"A5", -- 0x1FA0
    x"4E",x"85",x"38",x"E6",x"38",x"A9",x"01",x"C5", -- 0x1FA8
    x"37",x"F0",x"33",x"A4",x"49",x"30",x"0C",x"C4", -- 0x1FB0
    x"38",x"B0",x"2B",x"A9",x"00",x"85",x"49",x"C8", -- 0x1FB8
    x"98",x"D0",x"23",x"A5",x"37",x"C9",x"02",x"F0", -- 0x1FC0
    x"06",x"A9",x"01",x"C0",x"FF",x"D0",x"17",x"A9", -- 0x1FC8
    x"30",x"20",x"66",x"A0",x"A9",x"2E",x"20",x"66", -- 0x1FD0
    x"A0",x"A9",x"30",x"E6",x"49",x"F0",x"05",x"20", -- 0x1FD8
    x"66",x"A0",x"D0",x"F7",x"A9",x"80",x"85",x"4E", -- 0x1FE0
    x"20",x"40",x"A0",x"C6",x"4E",x"D0",x"05",x"A9", -- 0x1FE8
    x"2E",x"20",x"66",x"A0",x"C6",x"38",x"D0",x"F0", -- 0x1FF0
    x"A4",x"37",x"88",x"F0",x"18",x"88",x"F0",x"11", -- 0x1FF8
    x"A4",x"36",x"88",x"B9",x"00",x"06",x"C9",x"30", -- 0x2000
    x"F0",x"F8",x"C9",x"2E",x"F0",x"01",x"C8",x"84", -- 0x2008
    x"36",x"A5",x"49",x"F0",x"2A",x"A9",x"45",x"20", -- 0x2010
    x"66",x"A0",x"A5",x"49",x"10",x"0A",x"A9",x"2D", -- 0x2018
    x"20",x"66",x"A0",x"38",x"A9",x"00",x"E5",x"49", -- 0x2020
    x"20",x"52",x"A0",x"A5",x"37",x"F0",x"10",x"A9", -- 0x2028
    x"20",x"A4",x"49",x"30",x"03",x"20",x"66",x"A0", -- 0x2030
    x"E0",x"00",x"D0",x"03",x"4C",x"66",x"A0",x"60", -- 0x2038
    x"A5",x"31",x"4A",x"4A",x"4A",x"4A",x"20",x"64", -- 0x2040
    x"A0",x"A5",x"31",x"29",x"0F",x"85",x"31",x"4C", -- 0x2048
    x"97",x"A1",x"A2",x"FF",x"38",x"E8",x"E9",x"0A", -- 0x2050
    x"B0",x"FB",x"69",x"0A",x"48",x"8A",x"F0",x"03", -- 0x2058
    x"20",x"64",x"A0",x"68",x"09",x"30",x"86",x"3B", -- 0x2060
    x"A6",x"36",x"9D",x"00",x"06",x"A6",x"3B",x"E6", -- 0x2068
    x"36",x"60",x"18",x"86",x"35",x"20",x"DA",x"A1", -- 0x2070
    x"A9",x"FF",x"60",x"A2",x"00",x"86",x"31",x"86", -- 0x2078
    x"32",x"86",x"33",x"86",x"34",x"86",x"35",x"86", -- 0x2080
    x"48",x"86",x"49",x"C9",x"2E",x"F0",x"11",x"C9", -- 0x2088
    x"3A",x"B0",x"DF",x"E9",x"2F",x"30",x"DB",x"85", -- 0x2090
    x"35",x"C8",x"B1",x"19",x"C9",x"2E",x"D0",x"08", -- 0x2098
    x"A5",x"48",x"D0",x"44",x"E6",x"48",x"D0",x"F1", -- 0x20A0
    x"C9",x"45",x"F0",x"35",x"C9",x"3A",x"B0",x"38", -- 0x20A8
    x"E9",x"2F",x"90",x"34",x"A6",x"31",x"E0",x"18", -- 0x20B0
    x"90",x"08",x"A6",x"48",x"D0",x"DB",x"E6",x"49", -- 0x20B8
    x"B0",x"D7",x"A6",x"48",x"F0",x"02",x"C6",x"49", -- 0x20C0
    x"20",x"97",x"A1",x"65",x"35",x"85",x"35",x"90", -- 0x20C8
    x"C8",x"E6",x"34",x"D0",x"C4",x"E6",x"33",x"D0", -- 0x20D0
    x"C0",x"E6",x"32",x"D0",x"BC",x"E6",x"31",x"D0", -- 0x20D8
    x"B8",x"20",x"40",x"A1",x"65",x"49",x"85",x"49", -- 0x20E0
    x"84",x"1B",x"A5",x"49",x"05",x"48",x"F0",x"2F", -- 0x20E8
    x"20",x"DA",x"A1",x"F0",x"26",x"A9",x"A8",x"85", -- 0x20F0
    x"30",x"A9",x"00",x"85",x"2F",x"85",x"2E",x"20", -- 0x20F8
    x"03",x"A3",x"A5",x"49",x"30",x"0B",x"F0",x"10", -- 0x2100
    x"20",x"F4",x"A1",x"C6",x"49",x"D0",x"F9",x"F0", -- 0x2108
    x"07",x"20",x"4D",x"A2",x"E6",x"49",x"D0",x"F9", -- 0x2110
    x"20",x"5C",x"A6",x"38",x"A9",x"FF",x"60",x"A5", -- 0x2118
    x"32",x"85",x"2D",x"29",x"80",x"05",x"31",x"D0", -- 0x2120
    x"CC",x"A5",x"35",x"85",x"2A",x"A5",x"34",x"85", -- 0x2128
    x"2B",x"A5",x"33",x"85",x"2C",x"A9",x"40",x"38", -- 0x2130
    x"60",x"20",x"4B",x"A1",x"49",x"FF",x"38",x"60", -- 0x2138
    x"C8",x"B1",x"19",x"C9",x"2D",x"F0",x"F2",x"C9", -- 0x2140
    x"2B",x"D0",x"03",x"C8",x"B1",x"19",x"C9",x"3A", -- 0x2148
    x"B0",x"22",x"E9",x"2F",x"90",x"1E",x"85",x"4A", -- 0x2150
    x"C8",x"B1",x"19",x"C9",x"3A",x"B0",x"11",x"E9", -- 0x2158
    x"2F",x"90",x"0D",x"C8",x"85",x"43",x"A5",x"4A", -- 0x2160
    x"0A",x"0A",x"65",x"4A",x"0A",x"65",x"43",x"60", -- 0x2168
    x"A5",x"4A",x"18",x"60",x"A9",x"00",x"18",x"60", -- 0x2170
    x"A5",x"35",x"65",x"42",x"85",x"35",x"A5",x"34", -- 0x2178
    x"65",x"41",x"85",x"34",x"A5",x"33",x"65",x"40", -- 0x2180
    x"85",x"33",x"A5",x"32",x"65",x"3F",x"85",x"32", -- 0x2188
    x"A5",x"31",x"65",x"3E",x"85",x"31",x"60",x"48", -- 0x2190
    x"A6",x"34",x"A5",x"31",x"48",x"A5",x"32",x"48", -- 0x2198
    x"A5",x"33",x"48",x"A5",x"35",x"0A",x"26",x"34", -- 0x21A0
    x"26",x"33",x"26",x"32",x"26",x"31",x"0A",x"26", -- 0x21A8
    x"34",x"26",x"33",x"26",x"32",x"26",x"31",x"65", -- 0x21B0
    x"35",x"85",x"35",x"8A",x"65",x"34",x"85",x"34", -- 0x21B8
    x"68",x"65",x"33",x"85",x"33",x"68",x"65",x"32", -- 0x21C0
    x"85",x"32",x"68",x"65",x"31",x"06",x"35",x"26", -- 0x21C8
    x"34",x"26",x"33",x"26",x"32",x"2A",x"85",x"31", -- 0x21D0
    x"68",x"60",x"A5",x"31",x"05",x"32",x"05",x"33", -- 0x21D8
    x"05",x"34",x"05",x"35",x"F0",x"07",x"A5",x"2E", -- 0x21E0
    x"D0",x"09",x"A9",x"01",x"60",x"85",x"2E",x"85", -- 0x21E8
    x"30",x"85",x"2F",x"60",x"18",x"A5",x"30",x"69", -- 0x21F0
    x"03",x"85",x"30",x"90",x"02",x"E6",x"2F",x"20", -- 0x21F8
    x"1E",x"A2",x"20",x"42",x"A2",x"20",x"42",x"A2", -- 0x2200
    x"20",x"78",x"A1",x"90",x"10",x"66",x"31",x"66", -- 0x2208
    x"32",x"66",x"33",x"66",x"34",x"66",x"35",x"E6", -- 0x2210
    x"30",x"D0",x"02",x"E6",x"2F",x"60",x"A5",x"2E", -- 0x2218
    x"85",x"3B",x"A5",x"2F",x"85",x"3C",x"A5",x"30", -- 0x2220
    x"85",x"3D",x"A5",x"31",x"85",x"3E",x"A5",x"32", -- 0x2228
    x"85",x"3F",x"A5",x"33",x"85",x"40",x"A5",x"34", -- 0x2230
    x"85",x"41",x"A5",x"35",x"85",x"42",x"60",x"20", -- 0x2238
    x"1E",x"A2",x"46",x"3E",x"66",x"3F",x"66",x"40", -- 0x2240
    x"66",x"41",x"66",x"42",x"60",x"38",x"A5",x"30", -- 0x2248
    x"E9",x"04",x"85",x"30",x"B0",x"02",x"C6",x"2F", -- 0x2250
    x"20",x"3F",x"A2",x"20",x"08",x"A2",x"20",x"3F", -- 0x2258
    x"A2",x"20",x"42",x"A2",x"20",x"42",x"A2",x"20", -- 0x2260
    x"42",x"A2",x"20",x"08",x"A2",x"A9",x"00",x"85", -- 0x2268
    x"3E",x"A5",x"31",x"85",x"3F",x"A5",x"32",x"85", -- 0x2270
    x"40",x"A5",x"33",x"85",x"41",x"A5",x"34",x"85", -- 0x2278
    x"42",x"A5",x"35",x"2A",x"20",x"08",x"A2",x"A9", -- 0x2280
    x"00",x"85",x"3E",x"85",x"3F",x"A5",x"31",x"85", -- 0x2288
    x"40",x"A5",x"32",x"85",x"41",x"A5",x"33",x"85", -- 0x2290
    x"42",x"A5",x"34",x"2A",x"20",x"08",x"A2",x"A5", -- 0x2298
    x"32",x"2A",x"A5",x"31",x"65",x"35",x"85",x"35", -- 0x22A0
    x"90",x"13",x"E6",x"34",x"D0",x"0F",x"E6",x"33", -- 0x22A8
    x"D0",x"0B",x"E6",x"32",x"D0",x"07",x"E6",x"31", -- 0x22B0
    x"D0",x"03",x"4C",x"0B",x"A2",x"60",x"A2",x"00", -- 0x22B8
    x"86",x"35",x"86",x"2F",x"A5",x"2D",x"10",x"05", -- 0x22C0
    x"20",x"93",x"AD",x"A2",x"FF",x"86",x"2E",x"A5", -- 0x22C8
    x"2A",x"85",x"34",x"A5",x"2B",x"85",x"33",x"A5", -- 0x22D0
    x"2C",x"85",x"32",x"A5",x"2D",x"85",x"31",x"A9", -- 0x22D8
    x"A0",x"85",x"30",x"4C",x"03",x"A3",x"85",x"2E", -- 0x22E0
    x"85",x"30",x"85",x"2F",x"60",x"48",x"20",x"86", -- 0x22E8
    x"A6",x"68",x"F0",x"F8",x"10",x"07",x"85",x"2E", -- 0x22F0
    x"A9",x"00",x"38",x"E5",x"2E",x"85",x"31",x"A9", -- 0x22F8
    x"88",x"85",x"30",x"A5",x"31",x"30",x"E5",x"05", -- 0x2300
    x"32",x"05",x"33",x"05",x"34",x"05",x"35",x"F0", -- 0x2308
    x"D5",x"A5",x"30",x"A4",x"31",x"30",x"D5",x"D0", -- 0x2310
    x"21",x"A6",x"32",x"86",x"31",x"A6",x"33",x"86", -- 0x2318
    x"32",x"A6",x"34",x"86",x"33",x"A6",x"35",x"86", -- 0x2320
    x"34",x"84",x"35",x"38",x"E9",x"08",x"85",x"30", -- 0x2328
    x"B0",x"E1",x"C6",x"2F",x"90",x"DD",x"A4",x"31", -- 0x2330
    x"30",x"B2",x"06",x"35",x"26",x"34",x"26",x"33", -- 0x2338
    x"26",x"32",x"26",x"31",x"E9",x"00",x"85",x"30", -- 0x2340
    x"B0",x"EC",x"C6",x"2F",x"90",x"E8",x"A0",x"04", -- 0x2348
    x"B1",x"4B",x"85",x"41",x"88",x"B1",x"4B",x"85", -- 0x2350
    x"40",x"88",x"B1",x"4B",x"85",x"3F",x"88",x"B1", -- 0x2358
    x"4B",x"85",x"3B",x"88",x"84",x"42",x"84",x"3C", -- 0x2360
    x"B1",x"4B",x"85",x"3D",x"05",x"3B",x"05",x"3F", -- 0x2368
    x"05",x"40",x"05",x"41",x"F0",x"04",x"A5",x"3B", -- 0x2370
    x"09",x"80",x"85",x"3E",x"60",x"A9",x"71",x"D0", -- 0x2378
    x"06",x"A9",x"76",x"D0",x"02",x"A9",x"6C",x"85", -- 0x2380
    x"4B",x"A9",x"04",x"85",x"4C",x"A0",x"00",x"A5", -- 0x2388
    x"30",x"91",x"4B",x"C8",x"A5",x"2E",x"29",x"80", -- 0x2390
    x"85",x"2E",x"A5",x"31",x"29",x"7F",x"05",x"2E", -- 0x2398
    x"91",x"4B",x"A5",x"32",x"C8",x"91",x"4B",x"A5", -- 0x23A0
    x"33",x"C8",x"91",x"4B",x"A5",x"34",x"C8",x"91", -- 0x23A8
    x"4B",x"60",x"20",x"F5",x"A7",x"A0",x"04",x"B1", -- 0x23B0
    x"4B",x"85",x"34",x"88",x"B1",x"4B",x"85",x"33", -- 0x23B8
    x"88",x"B1",x"4B",x"85",x"32",x"88",x"B1",x"4B", -- 0x23C0
    x"85",x"2E",x"88",x"B1",x"4B",x"85",x"30",x"84", -- 0x23C8
    x"35",x"84",x"2F",x"05",x"2E",x"05",x"32",x"05", -- 0x23D0
    x"33",x"05",x"34",x"F0",x"04",x"A5",x"2E",x"09", -- 0x23D8
    x"80",x"85",x"31",x"60",x"20",x"FE",x"A3",x"A5", -- 0x23E0
    x"31",x"85",x"2D",x"A5",x"32",x"85",x"2C",x"A5", -- 0x23E8
    x"33",x"85",x"2B",x"A5",x"34",x"85",x"2A",x"60", -- 0x23F0
    x"20",x"1E",x"A2",x"4C",x"86",x"A6",x"A5",x"30", -- 0x23F8
    x"10",x"F6",x"20",x"53",x"A4",x"20",x"DA",x"A1", -- 0x2400
    x"D0",x"32",x"F0",x"5C",x"A5",x"30",x"C9",x"A0", -- 0x2408
    x"B0",x"54",x"C9",x"99",x"B0",x"26",x"69",x"08", -- 0x2410
    x"85",x"30",x"A5",x"40",x"85",x"41",x"A5",x"3F", -- 0x2418
    x"85",x"40",x"A5",x"3E",x"85",x"3F",x"A5",x"34", -- 0x2420
    x"85",x"3E",x"A5",x"33",x"85",x"34",x"A5",x"32", -- 0x2428
    x"85",x"33",x"A5",x"31",x"85",x"32",x"A9",x"00", -- 0x2430
    x"85",x"31",x"F0",x"D0",x"46",x"31",x"66",x"32", -- 0x2438
    x"66",x"33",x"66",x"34",x"66",x"3E",x"66",x"3F", -- 0x2440
    x"66",x"40",x"66",x"41",x"E6",x"30",x"D0",x"BC", -- 0x2448
    x"4C",x"6C",x"A6",x"A9",x"00",x"85",x"3B",x"85", -- 0x2450
    x"3C",x"85",x"3D",x"85",x"3E",x"85",x"3F",x"85", -- 0x2458
    x"40",x"85",x"41",x"85",x"42",x"60",x"D0",x"E8", -- 0x2460
    x"A5",x"2E",x"10",x"19",x"38",x"A9",x"00",x"E5", -- 0x2468
    x"34",x"85",x"34",x"A9",x"00",x"E5",x"33",x"85", -- 0x2470
    x"33",x"A9",x"00",x"E5",x"32",x"85",x"32",x"A9", -- 0x2478
    x"00",x"E5",x"31",x"85",x"31",x"60",x"A5",x"30", -- 0x2480
    x"30",x"07",x"A9",x"00",x"85",x"4A",x"4C",x"DA", -- 0x2488
    x"A1",x"20",x"FE",x"A3",x"A5",x"34",x"85",x"4A", -- 0x2490
    x"20",x"E8",x"A4",x"A9",x"80",x"85",x"30",x"A6", -- 0x2498
    x"31",x"10",x"10",x"45",x"2E",x"85",x"2E",x"10", -- 0x24A0
    x"05",x"E6",x"4A",x"4C",x"B0",x"A4",x"C6",x"4A", -- 0x24A8
    x"20",x"6C",x"A4",x"4C",x"03",x"A3",x"E6",x"34", -- 0x24B0
    x"D0",x"0C",x"E6",x"33",x"D0",x"08",x"E6",x"32", -- 0x24B8
    x"D0",x"04",x"E6",x"31",x"F0",x"8A",x"60",x"20", -- 0x24C0
    x"6C",x"A4",x"20",x"B6",x"A4",x"4C",x"6C",x"A4", -- 0x24C8
    x"20",x"FD",x"A4",x"4C",x"7E",x"AD",x"20",x"4E", -- 0x24D0
    x"A3",x"20",x"8D",x"A3",x"A5",x"3B",x"85",x"2E", -- 0x24D8
    x"A5",x"3C",x"85",x"2F",x"A5",x"3D",x"85",x"30", -- 0x24E0
    x"A5",x"3E",x"85",x"31",x"A5",x"3F",x"85",x"32", -- 0x24E8
    x"A5",x"40",x"85",x"33",x"A5",x"41",x"85",x"34", -- 0x24F0
    x"A5",x"42",x"85",x"35",x"60",x"20",x"7E",x"AD", -- 0x24F8
    x"20",x"4E",x"A3",x"F0",x"F7",x"20",x"0B",x"A5", -- 0x2500
    x"4C",x"5C",x"A6",x"20",x"DA",x"A1",x"F0",x"CC", -- 0x2508
    x"A0",x"00",x"38",x"A5",x"30",x"E5",x"3D",x"F0", -- 0x2510
    x"77",x"90",x"37",x"C9",x"25",x"B0",x"DD",x"48", -- 0x2518
    x"29",x"38",x"F0",x"19",x"4A",x"4A",x"4A",x"AA", -- 0x2520
    x"A5",x"41",x"85",x"42",x"A5",x"40",x"85",x"41", -- 0x2528
    x"A5",x"3F",x"85",x"40",x"A5",x"3E",x"85",x"3F", -- 0x2530
    x"84",x"3E",x"CA",x"D0",x"EB",x"68",x"29",x"07", -- 0x2538
    x"F0",x"4E",x"AA",x"46",x"3E",x"66",x"3F",x"66", -- 0x2540
    x"40",x"66",x"41",x"66",x"42",x"CA",x"D0",x"F3", -- 0x2548
    x"F0",x"3E",x"38",x"A5",x"3D",x"E5",x"30",x"C9", -- 0x2550
    x"25",x"B0",x"81",x"48",x"29",x"38",x"F0",x"19", -- 0x2558
    x"4A",x"4A",x"4A",x"AA",x"A5",x"34",x"85",x"35", -- 0x2560
    x"A5",x"33",x"85",x"34",x"A5",x"32",x"85",x"33", -- 0x2568
    x"A5",x"31",x"85",x"32",x"84",x"31",x"CA",x"D0", -- 0x2570
    x"EB",x"68",x"29",x"07",x"F0",x"0E",x"AA",x"46", -- 0x2578
    x"31",x"66",x"32",x"66",x"33",x"66",x"34",x"66", -- 0x2580
    x"35",x"CA",x"D0",x"F3",x"A5",x"3D",x"85",x"30", -- 0x2588
    x"A5",x"2E",x"45",x"3B",x"10",x"49",x"A5",x"31", -- 0x2590
    x"C5",x"3E",x"D0",x"1B",x"A5",x"32",x"C5",x"3F", -- 0x2598
    x"D0",x"15",x"A5",x"33",x"C5",x"40",x"D0",x"0F", -- 0x25A0
    x"A5",x"34",x"C5",x"41",x"D0",x"09",x"A5",x"35", -- 0x25A8
    x"C5",x"42",x"D0",x"03",x"4C",x"86",x"A6",x"B0", -- 0x25B0
    x"2A",x"38",x"A5",x"42",x"E5",x"35",x"85",x"35", -- 0x25B8
    x"A5",x"41",x"E5",x"34",x"85",x"34",x"A5",x"40", -- 0x25C0
    x"E5",x"33",x"85",x"33",x"A5",x"3F",x"E5",x"32", -- 0x25C8
    x"85",x"32",x"A5",x"3E",x"E5",x"31",x"85",x"31", -- 0x25D0
    x"A5",x"3B",x"85",x"2E",x"4C",x"03",x"A3",x"18", -- 0x25D8
    x"4C",x"08",x"A2",x"38",x"A5",x"35",x"E5",x"42", -- 0x25E0
    x"85",x"35",x"A5",x"34",x"E5",x"41",x"85",x"34", -- 0x25E8
    x"A5",x"33",x"E5",x"40",x"85",x"33",x"A5",x"32", -- 0x25F0
    x"E5",x"3F",x"85",x"32",x"A5",x"31",x"E5",x"3E", -- 0x25F8
    x"85",x"31",x"4C",x"03",x"A3",x"60",x"20",x"DA", -- 0x2600
    x"A1",x"F0",x"FA",x"20",x"4E",x"A3",x"D0",x"03", -- 0x2608
    x"4C",x"86",x"A6",x"18",x"A5",x"30",x"65",x"3D", -- 0x2610
    x"90",x"03",x"E6",x"2F",x"18",x"E9",x"7F",x"85", -- 0x2618
    x"30",x"B0",x"02",x"C6",x"2F",x"A2",x"05",x"A0", -- 0x2620
    x"00",x"B5",x"30",x"95",x"42",x"94",x"30",x"CA", -- 0x2628
    x"D0",x"F7",x"A5",x"2E",x"45",x"3B",x"85",x"2E", -- 0x2630
    x"A0",x"20",x"46",x"3E",x"66",x"3F",x"66",x"40", -- 0x2638
    x"66",x"41",x"66",x"42",x"06",x"46",x"26",x"45", -- 0x2640
    x"26",x"44",x"26",x"43",x"90",x"04",x"18",x"20", -- 0x2648
    x"78",x"A1",x"88",x"D0",x"E5",x"60",x"20",x"06", -- 0x2650
    x"A6",x"20",x"03",x"A3",x"A5",x"35",x"C9",x"80", -- 0x2658
    x"90",x"1A",x"F0",x"12",x"A9",x"FF",x"20",x"A4", -- 0x2660
    x"A2",x"4C",x"7C",x"A6",x"00",x"14",x"54",x"6F", -- 0x2668
    x"6F",x"20",x"62",x"69",x"67",x"00",x"A5",x"34", -- 0x2670
    x"09",x"01",x"85",x"34",x"A9",x"00",x"85",x"35", -- 0x2678
    x"A5",x"2F",x"F0",x"14",x"10",x"E6",x"A9",x"00", -- 0x2680
    x"85",x"2E",x"85",x"2F",x"85",x"30",x"85",x"31", -- 0x2688
    x"85",x"32",x"85",x"33",x"85",x"34",x"85",x"35", -- 0x2690
    x"60",x"20",x"86",x"A6",x"A0",x"80",x"84",x"31", -- 0x2698
    x"C8",x"84",x"30",x"98",x"60",x"20",x"85",x"A3", -- 0x26A0
    x"20",x"99",x"A6",x"D0",x"3A",x"20",x"DA",x"A1", -- 0x26A8
    x"F0",x"09",x"20",x"1E",x"A2",x"20",x"B5",x"A3", -- 0x26B0
    x"D0",x"37",x"60",x"4C",x"A7",x"99",x"20",x"FA", -- 0x26B8
    x"92",x"20",x"D3",x"A9",x"A5",x"4A",x"48",x"20", -- 0x26C0
    x"E9",x"A7",x"20",x"8D",x"A3",x"E6",x"4A",x"20", -- 0x26C8
    x"9E",x"A9",x"20",x"E9",x"A7",x"20",x"D6",x"A4", -- 0x26D0
    x"68",x"85",x"4A",x"20",x"9E",x"A9",x"20",x"E9", -- 0x26D8
    x"A7",x"20",x"E7",x"A6",x"A9",x"FF",x"60",x"20", -- 0x26E0
    x"DA",x"A1",x"F0",x"AC",x"20",x"4E",x"A3",x"F0", -- 0x26E8
    x"CA",x"A5",x"2E",x"45",x"3B",x"85",x"2E",x"38", -- 0x26F0
    x"A5",x"30",x"E5",x"3D",x"B0",x"03",x"C6",x"2F", -- 0x26F8
    x"38",x"69",x"80",x"85",x"30",x"90",x"03",x"E6", -- 0x2700
    x"2F",x"18",x"A2",x"20",x"B0",x"18",x"A5",x"31", -- 0x2708
    x"C5",x"3E",x"D0",x"10",x"A5",x"32",x"C5",x"3F", -- 0x2710
    x"D0",x"0A",x"A5",x"33",x"C5",x"40",x"D0",x"04", -- 0x2718
    x"A5",x"34",x"C5",x"41",x"90",x"19",x"A5",x"34", -- 0x2720
    x"E5",x"41",x"85",x"34",x"A5",x"33",x"E5",x"40", -- 0x2728
    x"85",x"33",x"A5",x"32",x"E5",x"3F",x"85",x"32", -- 0x2730
    x"A5",x"31",x"E5",x"3E",x"85",x"31",x"38",x"26", -- 0x2738
    x"46",x"26",x"45",x"26",x"44",x"26",x"43",x"06", -- 0x2740
    x"34",x"26",x"33",x"26",x"32",x"26",x"31",x"CA", -- 0x2748
    x"D0",x"BA",x"A2",x"07",x"B0",x"18",x"A5",x"31", -- 0x2750
    x"C5",x"3E",x"D0",x"10",x"A5",x"32",x"C5",x"3F", -- 0x2758
    x"D0",x"0A",x"A5",x"33",x"C5",x"40",x"D0",x"04", -- 0x2760
    x"A5",x"34",x"C5",x"41",x"90",x"19",x"A5",x"34", -- 0x2768
    x"E5",x"41",x"85",x"34",x"A5",x"33",x"E5",x"40", -- 0x2770
    x"85",x"33",x"A5",x"32",x"E5",x"3F",x"85",x"32", -- 0x2778
    x"A5",x"31",x"E5",x"3E",x"85",x"31",x"38",x"26", -- 0x2780
    x"35",x"06",x"34",x"26",x"33",x"26",x"32",x"26", -- 0x2788
    x"31",x"CA",x"D0",x"C0",x"06",x"35",x"A5",x"46", -- 0x2790
    x"85",x"34",x"A5",x"45",x"85",x"33",x"A5",x"44", -- 0x2798
    x"85",x"32",x"A5",x"43",x"85",x"31",x"4C",x"59", -- 0x27A0
    x"A6",x"00",x"15",x"2D",x"76",x"65",x"20",x"72", -- 0x27A8
    x"6F",x"6F",x"74",x"00",x"20",x"FA",x"92",x"20", -- 0x27B0
    x"DA",x"A1",x"F0",x"2A",x"30",x"EB",x"20",x"85", -- 0x27B8
    x"A3",x"A5",x"30",x"4A",x"69",x"40",x"85",x"30", -- 0x27C0
    x"A9",x"05",x"85",x"4A",x"20",x"ED",x"A7",x"20", -- 0x27C8
    x"8D",x"A3",x"A9",x"6C",x"85",x"4B",x"20",x"AD", -- 0x27D0
    x"A6",x"A9",x"71",x"85",x"4B",x"20",x"00",x"A5", -- 0x27D8
    x"C6",x"30",x"C6",x"4A",x"D0",x"E9",x"A9",x"FF", -- 0x27E0
    x"60",x"A9",x"7B",x"D0",x"0A",x"A9",x"71",x"D0", -- 0x27E8
    x"06",x"A9",x"76",x"D0",x"02",x"A9",x"6C",x"85", -- 0x27F0
    x"4B",x"A9",x"04",x"85",x"4C",x"60",x"20",x"FA", -- 0x27F8
    x"92",x"20",x"DA",x"A1",x"F0",x"02",x"10",x"0C", -- 0x2800
    x"00",x"16",x"4C",x"6F",x"67",x"20",x"72",x"61", -- 0x2808
    x"6E",x"67",x"65",x"00",x"20",x"53",x"A4",x"A0", -- 0x2810
    x"80",x"84",x"3B",x"84",x"3E",x"C8",x"84",x"3D", -- 0x2818
    x"A6",x"30",x"F0",x"06",x"A5",x"31",x"C9",x"B5", -- 0x2820
    x"90",x"02",x"E8",x"88",x"8A",x"48",x"84",x"30", -- 0x2828
    x"20",x"05",x"A5",x"A9",x"7B",x"20",x"87",x"A3", -- 0x2830
    x"A9",x"73",x"A0",x"A8",x"20",x"97",x"A8",x"20", -- 0x2838
    x"E9",x"A7",x"20",x"56",x"A6",x"20",x"56",x"A6", -- 0x2840
    x"20",x"00",x"A5",x"20",x"85",x"A3",x"68",x"38", -- 0x2848
    x"E9",x"81",x"20",x"ED",x"A2",x"A9",x"6E",x"85", -- 0x2850
    x"4B",x"A9",x"A8",x"85",x"4C",x"20",x"56",x"A6", -- 0x2858
    x"20",x"F5",x"A7",x"20",x"00",x"A5",x"A9",x"FF", -- 0x2860
    x"60",x"7F",x"5E",x"5B",x"D8",x"AA",x"80",x"31", -- 0x2868
    x"72",x"17",x"F8",x"06",x"7A",x"12",x"38",x"A5", -- 0x2870
    x"0B",x"88",x"79",x"0E",x"9F",x"F3",x"7C",x"2A", -- 0x2878
    x"AC",x"3F",x"B5",x"86",x"34",x"01",x"A2",x"7A", -- 0x2880
    x"7F",x"63",x"8E",x"37",x"EC",x"82",x"3F",x"FF", -- 0x2888
    x"FF",x"C1",x"7F",x"FF",x"FF",x"FF",x"FF",x"85", -- 0x2890
    x"4D",x"84",x"4E",x"20",x"85",x"A3",x"A0",x"00", -- 0x2898
    x"B1",x"4D",x"85",x"48",x"E6",x"4D",x"D0",x"02", -- 0x28A0
    x"E6",x"4E",x"A5",x"4D",x"85",x"4B",x"A5",x"4E", -- 0x28A8
    x"85",x"4C",x"20",x"B5",x"A3",x"20",x"F5",x"A7", -- 0x28B0
    x"20",x"AD",x"A6",x"18",x"A5",x"4D",x"69",x"05", -- 0x28B8
    x"85",x"4D",x"85",x"4B",x"A5",x"4E",x"69",x"00", -- 0x28C0
    x"85",x"4E",x"85",x"4C",x"20",x"00",x"A5",x"C6", -- 0x28C8
    x"48",x"D0",x"E2",x"60",x"20",x"DA",x"A8",x"4C", -- 0x28D0
    x"27",x"A9",x"20",x"FA",x"92",x"20",x"DA",x"A1", -- 0x28D8
    x"10",x"08",x"46",x"2E",x"20",x"EA",x"A8",x"4C", -- 0x28E0
    x"16",x"A9",x"20",x"81",x"A3",x"20",x"B1",x"A9", -- 0x28E8
    x"20",x"DA",x"A1",x"F0",x"09",x"20",x"F1",x"A7", -- 0x28F0
    x"20",x"AD",x"A6",x"4C",x"0A",x"A9",x"20",x"55", -- 0x28F8
    x"AA",x"20",x"B5",x"A3",x"A9",x"FF",x"60",x"20", -- 0x2900
    x"FA",x"92",x"20",x"DA",x"A1",x"F0",x"F5",x"10", -- 0x2908
    x"0A",x"46",x"2E",x"20",x"1B",x"A9",x"A9",x"80", -- 0x2910
    x"85",x"2E",x"60",x"A5",x"30",x"C9",x"81",x"90", -- 0x2918
    x"15",x"20",x"A5",x"A6",x"20",x"36",x"A9",x"20", -- 0x2920
    x"48",x"AA",x"20",x"00",x"A5",x"20",x"4C",x"AA", -- 0x2928
    x"20",x"00",x"A5",x"4C",x"7E",x"AD",x"A5",x"30", -- 0x2930
    x"C9",x"73",x"90",x"C8",x"20",x"81",x"A3",x"20", -- 0x2938
    x"53",x"A4",x"A9",x"80",x"85",x"3D",x"85",x"3E", -- 0x2940
    x"85",x"3B",x"20",x"05",x"A5",x"A9",x"5A",x"A0", -- 0x2948
    x"A9",x"20",x"97",x"A8",x"20",x"D1",x"AA",x"A9", -- 0x2950
    x"FF",x"60",x"09",x"85",x"A3",x"59",x"E8",x"67", -- 0x2958
    x"80",x"1C",x"9D",x"07",x"36",x"80",x"57",x"BB", -- 0x2960
    x"78",x"DF",x"80",x"CA",x"9A",x"0E",x"83",x"84", -- 0x2968
    x"8C",x"BB",x"CA",x"6E",x"81",x"95",x"96",x"06", -- 0x2970
    x"DE",x"81",x"0A",x"C7",x"6C",x"52",x"7F",x"7D", -- 0x2978
    x"AD",x"90",x"A1",x"82",x"FB",x"62",x"57",x"2F", -- 0x2980
    x"80",x"6D",x"63",x"38",x"2C",x"20",x"FA",x"92", -- 0x2988
    x"20",x"D3",x"A9",x"E6",x"4A",x"4C",x"9E",x"A9", -- 0x2990
    x"20",x"FA",x"92",x"20",x"D3",x"A9",x"A5",x"4A", -- 0x2998
    x"29",x"02",x"F0",x"06",x"20",x"AA",x"A9",x"4C", -- 0x29A0
    x"7E",x"AD",x"46",x"4A",x"90",x"15",x"20",x"C3", -- 0x29A8
    x"A9",x"20",x"85",x"A3",x"20",x"56",x"A6",x"20", -- 0x29B0
    x"8D",x"A3",x"20",x"99",x"A6",x"20",x"D0",x"A4", -- 0x29B8
    x"4C",x"B7",x"A7",x"20",x"81",x"A3",x"20",x"56", -- 0x29C0
    x"A6",x"A9",x"72",x"A0",x"AA",x"20",x"97",x"A8", -- 0x29C8
    x"4C",x"D1",x"AA",x"A5",x"30",x"C9",x"98",x"B0", -- 0x29D0
    x"5F",x"20",x"85",x"A3",x"20",x"55",x"AA",x"20", -- 0x29D8
    x"4E",x"A3",x"A5",x"2E",x"85",x"3B",x"C6",x"3D", -- 0x29E0
    x"20",x"05",x"A5",x"20",x"E7",x"A6",x"20",x"FE", -- 0x29E8
    x"A3",x"A5",x"34",x"85",x"4A",x"05",x"33",x"05", -- 0x29F0
    x"32",x"05",x"31",x"F0",x"38",x"A9",x"A0",x"85", -- 0x29F8
    x"30",x"A0",x"00",x"84",x"35",x"A5",x"31",x"85", -- 0x2A00
    x"2E",x"10",x"03",x"20",x"6C",x"A4",x"20",x"03", -- 0x2A08
    x"A3",x"20",x"7D",x"A3",x"20",x"48",x"AA",x"20", -- 0x2A10
    x"56",x"A6",x"20",x"F5",x"A7",x"20",x"00",x"A5", -- 0x2A18
    x"20",x"8D",x"A3",x"20",x"ED",x"A7",x"20",x"B5", -- 0x2A20
    x"A3",x"20",x"4C",x"AA",x"20",x"56",x"A6",x"20", -- 0x2A28
    x"F5",x"A7",x"4C",x"00",x"A5",x"4C",x"B2",x"A3", -- 0x2A30
    x"00",x"17",x"41",x"63",x"63",x"75",x"72",x"61", -- 0x2A38
    x"63",x"79",x"20",x"6C",x"6F",x"73",x"74",x"00", -- 0x2A40
    x"A9",x"59",x"D0",x"02",x"A9",x"5E",x"85",x"4B", -- 0x2A48
    x"A9",x"AA",x"85",x"4C",x"60",x"A9",x"63",x"D0", -- 0x2A50
    x"F5",x"81",x"C9",x"10",x"00",x"00",x"6F",x"15", -- 0x2A58
    x"77",x"7A",x"61",x"81",x"49",x"0F",x"DA",x"A2", -- 0x2A60
    x"7B",x"0E",x"FA",x"35",x"12",x"86",x"65",x"2E", -- 0x2A68
    x"E0",x"D3",x"05",x"84",x"8A",x"EA",x"0C",x"1B", -- 0x2A70
    x"84",x"1A",x"BE",x"BB",x"2B",x"84",x"37",x"45", -- 0x2A78
    x"55",x"AB",x"82",x"D5",x"55",x"57",x"7C",x"83", -- 0x2A80
    x"C0",x"00",x"00",x"05",x"81",x"00",x"00",x"00", -- 0x2A88
    x"00",x"20",x"FA",x"92",x"A5",x"30",x"C9",x"87", -- 0x2A90
    x"90",x"1E",x"D0",x"06",x"A4",x"31",x"C0",x"B3", -- 0x2A98
    x"90",x"16",x"A5",x"2E",x"10",x"06",x"20",x"86", -- 0x2AA0
    x"A6",x"A9",x"FF",x"60",x"00",x"18",x"45",x"78", -- 0x2AA8
    x"70",x"20",x"72",x"61",x"6E",x"67",x"65",x"00", -- 0x2AB0
    x"20",x"86",x"A4",x"20",x"DA",x"AA",x"20",x"81", -- 0x2AB8
    x"A3",x"A9",x"E4",x"85",x"4B",x"A9",x"AA",x"85", -- 0x2AC0
    x"4C",x"20",x"B5",x"A3",x"A5",x"4A",x"20",x"12", -- 0x2AC8
    x"AB",x"20",x"F1",x"A7",x"20",x"56",x"A6",x"A9", -- 0x2AD0
    x"FF",x"60",x"A9",x"E9",x"A0",x"AA",x"20",x"97", -- 0x2AD8
    x"A8",x"A9",x"FF",x"60",x"82",x"2D",x"F8",x"54", -- 0x2AE0
    x"58",x"07",x"83",x"E0",x"20",x"86",x"5B",x"82", -- 0x2AE8
    x"80",x"53",x"93",x"B8",x"83",x"20",x"00",x"06", -- 0x2AF0
    x"A1",x"82",x"00",x"00",x"21",x"63",x"82",x"C0", -- 0x2AF8
    x"00",x"00",x"02",x"82",x"80",x"00",x"00",x"0C", -- 0x2B00
    x"81",x"00",x"00",x"00",x"00",x"81",x"00",x"00", -- 0x2B08
    x"00",x"00",x"AA",x"10",x"09",x"CA",x"8A",x"49", -- 0x2B10
    x"FF",x"48",x"20",x"A5",x"A6",x"68",x"48",x"20", -- 0x2B18
    x"85",x"A3",x"20",x"99",x"A6",x"68",x"F0",x"0A", -- 0x2B20
    x"38",x"E9",x"01",x"48",x"20",x"56",x"A6",x"4C", -- 0x2B28
    x"25",x"AB",x"60",x"20",x"E3",x"92",x"A6",x"2A", -- 0x2B30
    x"A9",x"80",x"20",x"F4",x"FF",x"8A",x"4C",x"EA", -- 0x2B38
    x"AE",x"20",x"DD",x"92",x"20",x"94",x"BD",x"20", -- 0x2B40
    x"AE",x"8A",x"20",x"56",x"AE",x"20",x"F0",x"92", -- 0x2B48
    x"A5",x"2A",x"48",x"A5",x"2B",x"48",x"20",x"EA", -- 0x2B50
    x"BD",x"68",x"85",x"2D",x"68",x"85",x"2C",x"A2", -- 0x2B58
    x"2A",x"A9",x"09",x"20",x"F1",x"FF",x"A5",x"2E", -- 0x2B60
    x"30",x"33",x"4C",x"D8",x"AE",x"A9",x"86",x"20", -- 0x2B68
    x"F4",x"FF",x"8A",x"4C",x"D8",x"AE",x"A9",x"86", -- 0x2B70
    x"20",x"F4",x"FF",x"98",x"4C",x"D8",x"AE",x"20", -- 0x2B78
    x"DA",x"A1",x"F0",x"1E",x"10",x"1A",x"30",x"15", -- 0x2B80
    x"20",x"EC",x"AD",x"F0",x"59",x"30",x"F0",x"A5", -- 0x2B88
    x"2D",x"05",x"2C",x"05",x"2B",x"05",x"2A",x"F0", -- 0x2B90
    x"0C",x"A5",x"2D",x"10",x"03",x"4C",x"C4",x"AC", -- 0x2B98
    x"A9",x"01",x"4C",x"D8",x"AE",x"A9",x"40",x"60", -- 0x2BA0
    x"20",x"FE",x"A7",x"A0",x"69",x"A9",x"A8",x"D0", -- 0x2BA8
    x"07",x"20",x"FA",x"92",x"A0",x"68",x"A9",x"AA", -- 0x2BB0
    x"84",x"4B",x"85",x"4C",x"20",x"56",x"A6",x"A9", -- 0x2BB8
    x"FF",x"60",x"20",x"FA",x"92",x"A0",x"6D",x"A9", -- 0x2BC0
    x"AA",x"D0",x"ED",x"20",x"FE",x"A8",x"E6",x"30", -- 0x2BC8
    x"A8",x"60",x"20",x"E3",x"92",x"20",x"1E",x"8F", -- 0x2BD0
    x"85",x"2A",x"86",x"2B",x"84",x"2C",x"08",x"68", -- 0x2BD8
    x"85",x"2D",x"D8",x"A9",x"40",x"60",x"4C",x"0E", -- 0x2BE0
    x"8C",x"20",x"EC",x"AD",x"D0",x"F8",x"E6",x"36", -- 0x2BE8
    x"A4",x"36",x"A9",x"0D",x"99",x"FF",x"05",x"20", -- 0x2BF0
    x"B2",x"BD",x"A5",x"19",x"48",x"A5",x"1A",x"48", -- 0x2BF8
    x"A5",x"1B",x"48",x"A4",x"04",x"A6",x"05",x"C8", -- 0x2C00
    x"84",x"19",x"84",x"37",x"D0",x"01",x"E8",x"86", -- 0x2C08
    x"1A",x"86",x"38",x"A0",x"FF",x"84",x"3B",x"C8", -- 0x2C10
    x"84",x"1B",x"20",x"55",x"89",x"20",x"29",x"9B", -- 0x2C18
    x"20",x"DC",x"BD",x"68",x"85",x"1B",x"68",x"85", -- 0x2C20
    x"1A",x"68",x"85",x"19",x"A5",x"27",x"60",x"20", -- 0x2C28
    x"EC",x"AD",x"D0",x"67",x"A4",x"36",x"A9",x"00", -- 0x2C30
    x"99",x"00",x"06",x"A5",x"19",x"48",x"A5",x"1A", -- 0x2C38
    x"48",x"A5",x"1B",x"48",x"A9",x"00",x"85",x"1B", -- 0x2C40
    x"A9",x"00",x"85",x"19",x"A9",x"06",x"85",x"1A", -- 0x2C48
    x"20",x"8C",x"8A",x"C9",x"2D",x"F0",x"0F",x"C9", -- 0x2C50
    x"2B",x"D0",x"03",x"20",x"8C",x"8A",x"C6",x"1B", -- 0x2C58
    x"20",x"7B",x"A0",x"4C",x"73",x"AC",x"20",x"8C", -- 0x2C60
    x"8A",x"C6",x"1B",x"20",x"7B",x"A0",x"90",x"03", -- 0x2C68
    x"20",x"8F",x"AD",x"85",x"27",x"4C",x"23",x"AC", -- 0x2C70
    x"20",x"EC",x"AD",x"F0",x"1E",x"10",x"1B",x"A5", -- 0x2C78
    x"2E",x"08",x"20",x"FE",x"A3",x"28",x"10",x"0D", -- 0x2C80
    x"A5",x"3E",x"05",x"3F",x"05",x"40",x"05",x"41", -- 0x2C88
    x"F0",x"03",x"20",x"C7",x"A4",x"20",x"E7",x"A3", -- 0x2C90
    x"A9",x"40",x"60",x"4C",x"0E",x"8C",x"20",x"EC", -- 0x2C98
    x"AD",x"D0",x"F8",x"A5",x"36",x"F0",x"1D",x"AD", -- 0x2CA0
    x"00",x"06",x"4C",x"D8",x"AE",x"20",x"AD",x"AF", -- 0x2CA8
    x"C0",x"00",x"D0",x"10",x"8A",x"4C",x"EA",x"AE", -- 0x2CB0
    x"20",x"B5",x"BF",x"AA",x"A9",x"7F",x"20",x"F4", -- 0x2CB8
    x"FF",x"8A",x"F0",x"E6",x"A9",x"FF",x"85",x"2A", -- 0x2CC0
    x"85",x"2B",x"85",x"2C",x"85",x"2D",x"A9",x"40", -- 0x2CC8
    x"60",x"20",x"E3",x"92",x"A2",x"03",x"B5",x"2A", -- 0x2CD0
    x"49",x"FF",x"95",x"2A",x"CA",x"10",x"F7",x"A9", -- 0x2CD8
    x"40",x"60",x"20",x"29",x"9B",x"D0",x"B4",x"E0", -- 0x2CE0
    x"2C",x"D0",x"18",x"E6",x"1B",x"20",x"B2",x"BD", -- 0x2CE8
    x"20",x"29",x"9B",x"D0",x"A6",x"A9",x"01",x"85", -- 0x2CF0
    x"2A",x"E6",x"1B",x"E0",x"29",x"F0",x"13",x"E0", -- 0x2CF8
    x"2C",x"F0",x"03",x"4C",x"A2",x"8A",x"20",x"B2", -- 0x2D00
    x"BD",x"20",x"56",x"AE",x"20",x"F0",x"92",x"20", -- 0x2D08
    x"CB",x"BD",x"A0",x"00",x"A6",x"2A",x"D0",x"02", -- 0x2D10
    x"A2",x"01",x"86",x"2A",x"8A",x"CA",x"86",x"2D", -- 0x2D18
    x"18",x"65",x"04",x"85",x"37",x"98",x"65",x"05", -- 0x2D20
    x"85",x"38",x"B1",x"04",x"38",x"E5",x"2D",x"90", -- 0x2D28
    x"21",x"E5",x"36",x"90",x"1D",x"69",x"00",x"85", -- 0x2D30
    x"2B",x"20",x"DC",x"BD",x"A0",x"00",x"A6",x"36", -- 0x2D38
    x"F0",x"0B",x"B1",x"37",x"D9",x"00",x"06",x"D0", -- 0x2D40
    x"10",x"C8",x"CA",x"D0",x"F5",x"A5",x"2A",x"4C", -- 0x2D48
    x"D8",x"AE",x"20",x"DC",x"BD",x"A9",x"00",x"F0", -- 0x2D50
    x"F6",x"E6",x"2A",x"C6",x"2B",x"F0",x"F6",x"E6", -- 0x2D58
    x"37",x"D0",x"D9",x"E6",x"38",x"D0",x"D5",x"4C", -- 0x2D60
    x"0E",x"8C",x"20",x"EC",x"AD",x"F0",x"F8",x"30", -- 0x2D68
    x"06",x"24",x"2D",x"30",x"1E",x"10",x"33",x"20", -- 0x2D70
    x"DA",x"A1",x"10",x"0D",x"30",x"05",x"20",x"DA", -- 0x2D78
    x"A1",x"F0",x"06",x"A5",x"2E",x"49",x"80",x"85", -- 0x2D80
    x"2E",x"A9",x"FF",x"60",x"20",x"02",x"AE",x"F0", -- 0x2D88
    x"D6",x"30",x"EB",x"38",x"A9",x"00",x"A8",x"E5", -- 0x2D90
    x"2A",x"85",x"2A",x"98",x"E5",x"2B",x"85",x"2B", -- 0x2D98
    x"98",x"E5",x"2C",x"85",x"2C",x"98",x"E5",x"2D", -- 0x2DA0
    x"85",x"2D",x"A9",x"40",x"60",x"20",x"8C",x"8A", -- 0x2DA8
    x"C9",x"22",x"F0",x"15",x"A2",x"00",x"B1",x"19", -- 0x2DB0
    x"9D",x"00",x"06",x"C8",x"E8",x"C9",x"0D",x"F0", -- 0x2DB8
    x"04",x"C9",x"2C",x"D0",x"F1",x"88",x"4C",x"E1", -- 0x2DC0
    x"AD",x"A2",x"00",x"C8",x"B1",x"19",x"C9",x"0D", -- 0x2DC8
    x"F0",x"17",x"C8",x"9D",x"00",x"06",x"E8",x"C9", -- 0x2DD0
    x"22",x"D0",x"F1",x"B1",x"19",x"C9",x"22",x"F0", -- 0x2DD8
    x"EA",x"CA",x"86",x"36",x"84",x"1B",x"A9",x"00", -- 0x2DE0
    x"60",x"4C",x"98",x"8E",x"A4",x"1B",x"E6",x"1B", -- 0x2DE8
    x"B1",x"19",x"C9",x"20",x"F0",x"F6",x"C9",x"2D", -- 0x2DF0
    x"F0",x"92",x"C9",x"22",x"F0",x"CB",x"C9",x"2B", -- 0x2DF8
    x"D0",x"03",x"20",x"8C",x"8A",x"C9",x"8E",x"90", -- 0x2E00
    x"07",x"C9",x"C6",x"B0",x"36",x"4C",x"B1",x"8B", -- 0x2E08
    x"C9",x"3F",x"B0",x"0C",x"C9",x"2E",x"B0",x"12", -- 0x2E10
    x"C9",x"26",x"F0",x"51",x"C9",x"28",x"F0",x"36", -- 0x2E18
    x"C6",x"1B",x"20",x"DD",x"95",x"F0",x"09",x"4C", -- 0x2E20
    x"2C",x"B3",x"20",x"7B",x"A0",x"90",x"14",x"60", -- 0x2E28
    x"A5",x"28",x"29",x"02",x"D0",x"0D",x"B0",x"0B", -- 0x2E30
    x"86",x"1B",x"AD",x"40",x"04",x"AC",x"41",x"04", -- 0x2E38
    x"4C",x"EA",x"AE",x"00",x"1A",x"4E",x"6F",x"20", -- 0x2E40
    x"73",x"75",x"63",x"68",x"20",x"76",x"61",x"72", -- 0x2E48
    x"69",x"61",x"62",x"6C",x"65",x"00",x"20",x"29", -- 0x2E50
    x"9B",x"E6",x"1B",x"E0",x"29",x"D0",x"02",x"A8", -- 0x2E58
    x"60",x"00",x"1B",x"4D",x"69",x"73",x"73",x"69", -- 0x2E60
    x"6E",x"67",x"20",x"29",x"00",x"A2",x"00",x"86", -- 0x2E68
    x"2A",x"86",x"2B",x"86",x"2C",x"86",x"2D",x"A4", -- 0x2E70
    x"1B",x"B1",x"19",x"C9",x"30",x"90",x"23",x"C9", -- 0x2E78
    x"3A",x"90",x"0A",x"E9",x"37",x"C9",x"0A",x"90", -- 0x2E80
    x"19",x"C9",x"10",x"B0",x"15",x"0A",x"0A",x"0A", -- 0x2E88
    x"0A",x"A2",x"03",x"0A",x"26",x"2A",x"26",x"2B", -- 0x2E90
    x"26",x"2C",x"26",x"2D",x"CA",x"10",x"F4",x"C8", -- 0x2E98
    x"D0",x"D7",x"8A",x"10",x"05",x"84",x"1B",x"A9", -- 0x2EA0
    x"40",x"60",x"00",x"1C",x"42",x"61",x"64",x"20", -- 0x2EA8
    x"48",x"45",x"58",x"00",x"A2",x"2A",x"A0",x"00", -- 0x2EB0
    x"A9",x"01",x"20",x"F1",x"FF",x"A9",x"40",x"60", -- 0x2EB8
    x"A9",x"00",x"A4",x"18",x"4C",x"EA",x"AE",x"4C", -- 0x2EC0
    x"43",x"AE",x"A9",x"00",x"F0",x"0A",x"4C",x"0E", -- 0x2EC8
    x"8C",x"20",x"EC",x"AD",x"D0",x"F8",x"A5",x"36", -- 0x2ED0
    x"A0",x"00",x"F0",x"0E",x"A4",x"1B",x"B1",x"19", -- 0x2ED8
    x"C9",x"50",x"D0",x"E3",x"E6",x"1B",x"A5",x"12", -- 0x2EE0
    x"A4",x"13",x"85",x"2A",x"84",x"2B",x"A9",x"00", -- 0x2EE8
    x"85",x"2C",x"85",x"2D",x"A9",x"40",x"60",x"A5", -- 0x2EF0
    x"1E",x"4C",x"D8",x"AE",x"A5",x"00",x"A4",x"01", -- 0x2EF8
    x"4C",x"EA",x"AE",x"A5",x"06",x"A4",x"07",x"4C", -- 0x2F00
    x"EA",x"AE",x"E6",x"1B",x"20",x"56",x"AE",x"20", -- 0x2F08
    x"F0",x"92",x"A5",x"2D",x"30",x"29",x"05",x"2C", -- 0x2F10
    x"05",x"2B",x"D0",x"08",x"A5",x"2A",x"F0",x"4C", -- 0x2F18
    x"C9",x"01",x"F0",x"45",x"20",x"BE",x"A2",x"20", -- 0x2F20
    x"51",x"BD",x"20",x"69",x"AF",x"20",x"7E",x"BD", -- 0x2F28
    x"20",x"06",x"A6",x"20",x"03",x"A3",x"20",x"E4", -- 0x2F30
    x"A3",x"20",x"22",x"92",x"A9",x"40",x"60",x"A2", -- 0x2F38
    x"0D",x"20",x"44",x"BE",x"A9",x"40",x"85",x"11", -- 0x2F40
    x"60",x"A4",x"1B",x"B1",x"19",x"C9",x"28",x"F0", -- 0x2F48
    x"B9",x"20",x"87",x"AF",x"A2",x"0D",x"B5",x"00", -- 0x2F50
    x"85",x"2A",x"B5",x"01",x"85",x"2B",x"B5",x"02", -- 0x2F58
    x"85",x"2C",x"B5",x"03",x"85",x"2D",x"A9",x"40", -- 0x2F60
    x"60",x"20",x"87",x"AF",x"A2",x"00",x"86",x"2E", -- 0x2F68
    x"86",x"2F",x"86",x"35",x"A9",x"80",x"85",x"30", -- 0x2F70
    x"B5",x"0D",x"95",x"31",x"E8",x"E0",x"04",x"D0", -- 0x2F78
    x"F7",x"20",x"59",x"A6",x"A9",x"FF",x"60",x"A0", -- 0x2F80
    x"20",x"A5",x"0F",x"4A",x"4A",x"4A",x"45",x"11", -- 0x2F88
    x"6A",x"26",x"0D",x"26",x"0E",x"26",x"0F",x"26", -- 0x2F90
    x"10",x"26",x"11",x"88",x"D0",x"EB",x"60",x"A4", -- 0x2F98
    x"09",x"A5",x"08",x"4C",x"EA",x"AE",x"A0",x"00", -- 0x2FA0
    x"B1",x"FD",x"4C",x"EA",x"AE",x"20",x"E3",x"92", -- 0x2FA8
    x"A9",x"81",x"A6",x"2A",x"A4",x"2B",x"4C",x"F4", -- 0x2FB0
    x"FF",x"20",x"E0",x"FF",x"4C",x"D8",x"AE",x"20", -- 0x2FB8
    x"E0",x"FF",x"8D",x"00",x"06",x"A9",x"01",x"85", -- 0x2FC0
    x"36",x"A9",x"00",x"60",x"20",x"29",x"9B",x"D0", -- 0x2FC8
    x"62",x"E0",x"2C",x"D0",x"61",x"E6",x"1B",x"20", -- 0x2FD0
    x"B2",x"BD",x"20",x"56",x"AE",x"20",x"F0",x"92", -- 0x2FD8
    x"20",x"CB",x"BD",x"A5",x"2A",x"C5",x"36",x"B0", -- 0x2FE0
    x"02",x"85",x"36",x"A9",x"00",x"60",x"20",x"29", -- 0x2FE8
    x"9B",x"D0",x"40",x"E0",x"2C",x"D0",x"3F",x"E6", -- 0x2FF0
    x"1B",x"20",x"B2",x"BD",x"20",x"56",x"AE",x"20", -- 0x2FF8
    x"F0",x"92",x"20",x"CB",x"BD",x"A5",x"36",x"38", -- 0x3000
    x"E5",x"2A",x"90",x"17",x"F0",x"17",x"AA",x"A5", -- 0x3008
    x"2A",x"85",x"36",x"F0",x"10",x"A0",x"00",x"BD", -- 0x3010
    x"00",x"06",x"99",x"00",x"06",x"E8",x"C8",x"C6", -- 0x3018
    x"2A",x"D0",x"F4",x"A9",x"00",x"60",x"20",x"AD", -- 0x3020
    x"AF",x"8A",x"C0",x"00",x"F0",x"94",x"A9",x"00", -- 0x3028
    x"85",x"36",x"60",x"4C",x"0E",x"8C",x"4C",x"A2", -- 0x3030
    x"8A",x"20",x"29",x"9B",x"D0",x"F5",x"E0",x"2C", -- 0x3038
    x"D0",x"F4",x"20",x"B2",x"BD",x"E6",x"1B",x"20", -- 0x3040
    x"DD",x"92",x"A5",x"2A",x"48",x"A9",x"FF",x"85", -- 0x3048
    x"2A",x"E6",x"1B",x"E0",x"29",x"F0",x"0A",x"E0", -- 0x3050
    x"2C",x"D0",x"DB",x"20",x"56",x"AE",x"20",x"F0", -- 0x3058
    x"92",x"20",x"CB",x"BD",x"68",x"A8",x"18",x"F0", -- 0x3060
    x"06",x"E5",x"36",x"B0",x"C1",x"88",x"98",x"85", -- 0x3068
    x"2C",x"AA",x"A0",x"00",x"A5",x"36",x"38",x"E5", -- 0x3070
    x"2C",x"C5",x"2A",x"B0",x"02",x"85",x"2A",x"A5", -- 0x3078
    x"2A",x"F0",x"AB",x"BD",x"00",x"06",x"99",x"00", -- 0x3080
    x"06",x"C8",x"E8",x"C4",x"2A",x"D0",x"F4",x"84", -- 0x3088
    x"36",x"A9",x"00",x"60",x"20",x"8C",x"8A",x"A0", -- 0x3090
    x"FF",x"C9",x"7E",x"F0",x"04",x"A0",x"00",x"C6", -- 0x3098
    x"1B",x"98",x"48",x"20",x"EC",x"AD",x"F0",x"17", -- 0x30A0
    x"A8",x"68",x"85",x"15",x"AD",x"03",x"04",x"D0", -- 0x30A8
    x"08",x"85",x"37",x"20",x"F9",x"9E",x"A9",x"00", -- 0x30B0
    x"60",x"20",x"DF",x"9E",x"A9",x"00",x"60",x"4C", -- 0x30B8
    x"0E",x"8C",x"20",x"DD",x"92",x"20",x"94",x"BD", -- 0x30C0
    x"20",x"AE",x"8A",x"20",x"56",x"AE",x"D0",x"EF", -- 0x30C8
    x"20",x"EA",x"BD",x"A4",x"36",x"F0",x"1E",x"A5", -- 0x30D0
    x"2A",x"F0",x"1D",x"C6",x"2A",x"F0",x"16",x"A2", -- 0x30D8
    x"00",x"BD",x"00",x"06",x"99",x"00",x"06",x"E8", -- 0x30E0
    x"C8",x"F0",x"10",x"E4",x"36",x"90",x"F2",x"C6", -- 0x30E8
    x"2A",x"D0",x"EC",x"84",x"36",x"A9",x"00",x"60", -- 0x30F0
    x"85",x"36",x"60",x"4C",x"03",x"9C",x"68",x"85", -- 0x30F8
    x"0C",x"68",x"85",x"0B",x"00",x"1D",x"4E",x"6F", -- 0x3100
    x"20",x"73",x"75",x"63",x"68",x"20",x"A4",x"2F", -- 0x3108
    x"F2",x"00",x"A5",x"18",x"85",x"0C",x"A9",x"00", -- 0x3110
    x"85",x"0B",x"A0",x"01",x"B1",x"0B",x"30",x"DE", -- 0x3118
    x"A0",x"03",x"C8",x"B1",x"0B",x"C9",x"20",x"F0", -- 0x3120
    x"F9",x"C9",x"DD",x"F0",x"0F",x"A0",x"03",x"B1", -- 0x3128
    x"0B",x"18",x"65",x"0B",x"85",x"0B",x"90",x"E2", -- 0x3130
    x"E6",x"0C",x"B0",x"DE",x"C8",x"84",x"0A",x"20", -- 0x3138
    x"97",x"8A",x"98",x"AA",x"18",x"65",x"0B",x"A4", -- 0x3140
    x"0C",x"90",x"02",x"C8",x"18",x"E9",x"00",x"85", -- 0x3148
    x"3C",x"98",x"E9",x"00",x"85",x"3D",x"A0",x"00", -- 0x3150
    x"C8",x"E8",x"B1",x"3C",x"D1",x"37",x"D0",x"CD", -- 0x3158
    x"C4",x"39",x"D0",x"F4",x"C8",x"B1",x"3C",x"20", -- 0x3160
    x"26",x"89",x"B0",x"C1",x"8A",x"A8",x"20",x"6D", -- 0x3168
    x"98",x"20",x"ED",x"94",x"A2",x"01",x"20",x"31", -- 0x3170
    x"95",x"A0",x"00",x"A5",x"0B",x"91",x"02",x"C8", -- 0x3178
    x"A5",x"0C",x"91",x"02",x"20",x"39",x"95",x"4C", -- 0x3180
    x"F4",x"B1",x"00",x"1E",x"42",x"61",x"64",x"20", -- 0x3188
    x"63",x"61",x"6C",x"6C",x"00",x"A9",x"A4",x"85", -- 0x3190
    x"27",x"BA",x"8A",x"18",x"65",x"04",x"20",x"2E", -- 0x3198
    x"BE",x"A0",x"00",x"8A",x"91",x"04",x"E8",x"C8", -- 0x31A0
    x"BD",x"00",x"01",x"91",x"04",x"E0",x"FF",x"D0", -- 0x31A8
    x"F5",x"9A",x"A5",x"27",x"48",x"A5",x"0A",x"48", -- 0x31B0
    x"A5",x"0B",x"48",x"A5",x"0C",x"48",x"A5",x"1B", -- 0x31B8
    x"AA",x"18",x"65",x"19",x"A4",x"1A",x"90",x"02", -- 0x31C0
    x"C8",x"18",x"E9",x"01",x"85",x"37",x"98",x"E9", -- 0x31C8
    x"00",x"85",x"38",x"A0",x"02",x"20",x"5B",x"95", -- 0x31D0
    x"C0",x"02",x"F0",x"AE",x"86",x"1B",x"88",x"84", -- 0x31D8
    x"39",x"20",x"5B",x"94",x"D0",x"03",x"4C",x"12", -- 0x31E0
    x"B1",x"A0",x"00",x"B1",x"2A",x"85",x"0B",x"C8", -- 0x31E8
    x"B1",x"2A",x"85",x"0C",x"A9",x"00",x"48",x"85", -- 0x31F0
    x"0A",x"20",x"97",x"8A",x"C9",x"28",x"F0",x"4D", -- 0x31F8
    x"C6",x"0A",x"A5",x"1B",x"48",x"A5",x"19",x"48", -- 0x3200
    x"A5",x"1A",x"48",x"20",x"A3",x"8B",x"68",x"85", -- 0x3208
    x"1A",x"68",x"85",x"19",x"68",x"85",x"1B",x"68", -- 0x3210
    x"F0",x"0C",x"85",x"3F",x"20",x"0B",x"BE",x"20", -- 0x3218
    x"C1",x"8C",x"C6",x"3F",x"D0",x"F6",x"68",x"85", -- 0x3220
    x"0C",x"68",x"85",x"0B",x"68",x"85",x"0A",x"68", -- 0x3228
    x"A0",x"00",x"B1",x"04",x"AA",x"9A",x"C8",x"E8", -- 0x3230
    x"B1",x"04",x"9D",x"00",x"01",x"E0",x"FF",x"D0", -- 0x3238
    x"F5",x"98",x"65",x"04",x"85",x"04",x"90",x"02", -- 0x3240
    x"E6",x"05",x"A5",x"27",x"60",x"A5",x"1B",x"48", -- 0x3248
    x"A5",x"19",x"48",x"A5",x"1A",x"48",x"20",x"82", -- 0x3250
    x"95",x"F0",x"5A",x"A5",x"1B",x"85",x"0A",x"68", -- 0x3258
    x"85",x"1A",x"68",x"85",x"19",x"68",x"85",x"1B", -- 0x3260
    x"68",x"AA",x"A5",x"2C",x"48",x"A5",x"2B",x"48", -- 0x3268
    x"A5",x"2A",x"48",x"E8",x"8A",x"48",x"20",x"0D", -- 0x3270
    x"B3",x"20",x"97",x"8A",x"C9",x"2C",x"F0",x"CD", -- 0x3278
    x"C9",x"29",x"D0",x"31",x"A9",x"00",x"48",x"20", -- 0x3280
    x"8C",x"8A",x"C9",x"28",x"D0",x"27",x"20",x"29", -- 0x3288
    x"9B",x"20",x"90",x"BD",x"A5",x"27",x"85",x"2D", -- 0x3290
    x"20",x"94",x"BD",x"68",x"AA",x"E8",x"8A",x"48", -- 0x3298
    x"20",x"8C",x"8A",x"C9",x"2C",x"F0",x"E7",x"C9", -- 0x32A0
    x"29",x"D0",x"0A",x"68",x"68",x"85",x"4D",x"85", -- 0x32A8
    x"4E",x"E4",x"4D",x"F0",x"15",x"A2",x"FB",x"9A", -- 0x32B0
    x"68",x"85",x"0C",x"68",x"85",x"0B",x"00",x"1F", -- 0x32B8
    x"41",x"72",x"67",x"75",x"6D",x"65",x"6E",x"74", -- 0x32C0
    x"73",x"00",x"20",x"EA",x"BD",x"68",x"85",x"2A", -- 0x32C8
    x"68",x"85",x"2B",x"68",x"85",x"2C",x"30",x"21", -- 0x32D0
    x"A5",x"2D",x"F0",x"D9",x"85",x"27",x"A2",x"37", -- 0x32D8
    x"20",x"44",x"BE",x"A5",x"27",x"10",x"09",x"20", -- 0x32E0
    x"7E",x"BD",x"20",x"B5",x"A3",x"4C",x"F3",x"B2", -- 0x32E8
    x"20",x"EA",x"BD",x"20",x"B7",x"B4",x"4C",x"03", -- 0x32F0
    x"B3",x"A5",x"2D",x"D0",x"B8",x"20",x"CB",x"BD", -- 0x32F8
    x"20",x"21",x"8C",x"C6",x"4D",x"D0",x"C3",x"A5", -- 0x3300
    x"4E",x"48",x"4C",x"02",x"B2",x"A4",x"2C",x"C0", -- 0x3308
    x"04",x"D0",x"05",x"A2",x"37",x"20",x"44",x"BE", -- 0x3310
    x"20",x"2C",x"B3",x"08",x"20",x"90",x"BD",x"28", -- 0x3318
    x"F0",x"07",x"30",x"05",x"A2",x"37",x"20",x"56", -- 0x3320
    x"AF",x"4C",x"94",x"BD",x"A4",x"2C",x"30",x"54", -- 0x3328
    x"F0",x"1D",x"C0",x"05",x"F0",x"1E",x"A0",x"03", -- 0x3330
    x"B1",x"2A",x"85",x"2D",x"88",x"B1",x"2A",x"85", -- 0x3338
    x"2C",x"88",x"B1",x"2A",x"AA",x"88",x"B1",x"2A", -- 0x3340
    x"85",x"2A",x"86",x"2B",x"A9",x"40",x"60",x"B1", -- 0x3348
    x"2A",x"4C",x"EA",x"AE",x"88",x"B1",x"2A",x"85", -- 0x3350
    x"34",x"88",x"B1",x"2A",x"85",x"33",x"88",x"B1", -- 0x3358
    x"2A",x"85",x"32",x"88",x"B1",x"2A",x"85",x"2E", -- 0x3360
    x"88",x"B1",x"2A",x"85",x"30",x"84",x"35",x"84", -- 0x3368
    x"2F",x"05",x"2E",x"05",x"32",x"05",x"33",x"05", -- 0x3370
    x"34",x"F0",x"04",x"A5",x"2E",x"09",x"80",x"85", -- 0x3378
    x"31",x"A9",x"FF",x"60",x"C0",x"80",x"F0",x"1F", -- 0x3380
    x"A0",x"03",x"B1",x"2A",x"85",x"36",x"F0",x"16", -- 0x3388
    x"A0",x"01",x"B1",x"2A",x"85",x"38",x"88",x"B1", -- 0x3390
    x"2A",x"85",x"37",x"A4",x"36",x"88",x"B1",x"37", -- 0x3398
    x"99",x"00",x"06",x"98",x"D0",x"F7",x"60",x"A5", -- 0x33A0
    x"2B",x"F0",x"15",x"A0",x"00",x"B1",x"2A",x"99", -- 0x33A8
    x"00",x"06",x"49",x"0D",x"F0",x"04",x"C8",x"D0", -- 0x33B0
    x"F4",x"98",x"84",x"36",x"60",x"20",x"E3",x"92", -- 0x33B8
    x"A5",x"2A",x"4C",x"C2",x"AF",x"A0",x"00",x"84", -- 0x33C0
    x"08",x"84",x"09",x"A6",x"18",x"86",x"38",x"84", -- 0x33C8
    x"37",x"A6",x"0C",x"E0",x"07",x"F0",x"2A",x"A6", -- 0x33D0
    x"0B",x"20",x"42",x"89",x"C9",x"0D",x"D0",x"19", -- 0x33D8
    x"E4",x"37",x"A5",x"0C",x"E5",x"38",x"90",x"19", -- 0x33E0
    x"20",x"42",x"89",x"09",x"00",x"30",x"12",x"85", -- 0x33E8
    x"09",x"20",x"42",x"89",x"85",x"08",x"20",x"42", -- 0x33F0
    x"89",x"E4",x"37",x"A5",x"0C",x"E5",x"38",x"B0", -- 0x33F8
    x"D8",x"60",x"20",x"C5",x"B3",x"84",x"20",x"B1", -- 0x3400
    x"FD",x"D0",x"08",x"A9",x"33",x"85",x"16",x"A9", -- 0x3408
    x"B4",x"85",x"17",x"A5",x"16",x"85",x"0B",x"A5", -- 0x3410
    x"17",x"85",x"0C",x"20",x"3A",x"BD",x"AA",x"86", -- 0x3418
    x"0A",x"A9",x"DA",x"20",x"F4",x"FF",x"A9",x"7E", -- 0x3420
    x"20",x"F4",x"FF",x"A2",x"FF",x"86",x"28",x"9A", -- 0x3428
    x"4C",x"A3",x"8B",x"F6",x"3A",x"E7",x"9E",x"F1", -- 0x3430
    x"22",x"20",x"61",x"74",x"20",x"6C",x"69",x"6E", -- 0x3438
    x"65",x"20",x"22",x"3B",x"9E",x"3A",x"E0",x"8B", -- 0x3440
    x"F1",x"3A",x"E0",x"0D",x"20",x"21",x"88",x"A2", -- 0x3448
    x"03",x"A5",x"2A",x"48",x"A5",x"2B",x"48",x"8A", -- 0x3450
    x"48",x"20",x"DA",x"92",x"68",x"AA",x"CA",x"D0", -- 0x3458
    x"F0",x"20",x"52",x"98",x"A5",x"2A",x"85",x"3D", -- 0x3460
    x"A5",x"2B",x"85",x"3E",x"A0",x"07",x"A2",x"05", -- 0x3468
    x"D0",x"1D",x"20",x"21",x"88",x"A2",x"0D",x"A5", -- 0x3470
    x"2A",x"48",x"8A",x"48",x"20",x"DA",x"92",x"68", -- 0x3478
    x"AA",x"CA",x"D0",x"F3",x"20",x"52",x"98",x"A5", -- 0x3480
    x"2A",x"85",x"44",x"A2",x"0C",x"A0",x"08",x"68", -- 0x3488
    x"95",x"37",x"CA",x"10",x"FA",x"98",x"A2",x"37", -- 0x3490
    x"A0",x"00",x"20",x"F1",x"FF",x"4C",x"9B",x"8B", -- 0x3498
    x"20",x"21",x"88",x"20",x"52",x"98",x"A4",x"2A", -- 0x34A0
    x"88",x"84",x"23",x"4C",x"9B",x"8B",x"4C",x"0E", -- 0x34A8
    x"8C",x"20",x"29",x"9B",x"20",x"0B",x"BE",x"A5", -- 0x34B0
    x"39",x"C9",x"05",x"F0",x"23",x"A5",x"27",x"F0", -- 0x34B8
    x"ED",x"10",x"03",x"20",x"E4",x"A3",x"A0",x"00", -- 0x34C0
    x"A5",x"2A",x"91",x"37",x"A5",x"39",x"F0",x"0F", -- 0x34C8
    x"A5",x"2B",x"C8",x"91",x"37",x"A5",x"2C",x"C8", -- 0x34D0
    x"91",x"37",x"A5",x"2D",x"C8",x"91",x"37",x"60", -- 0x34D8
    x"A5",x"27",x"F0",x"CA",x"30",x"03",x"20",x"BE", -- 0x34E0
    x"A2",x"A0",x"00",x"A5",x"30",x"91",x"37",x"C8", -- 0x34E8
    x"A5",x"2E",x"29",x"80",x"85",x"2E",x"A5",x"31", -- 0x34F0
    x"29",x"7F",x"05",x"2E",x"91",x"37",x"C8",x"A5", -- 0x34F8
    x"32",x"91",x"37",x"C8",x"A5",x"33",x"91",x"37", -- 0x3500
    x"C8",x"A5",x"34",x"91",x"37",x"60",x"85",x"37", -- 0x3508
    x"C9",x"80",x"90",x"44",x"A9",x"71",x"85",x"38", -- 0x3510
    x"A9",x"80",x"85",x"39",x"84",x"3A",x"A0",x"00", -- 0x3518
    x"C8",x"B1",x"38",x"10",x"FB",x"C5",x"37",x"F0", -- 0x3520
    x"0D",x"C8",x"98",x"38",x"65",x"38",x"85",x"38", -- 0x3528
    x"90",x"EC",x"E6",x"39",x"B0",x"E8",x"A0",x"00", -- 0x3530
    x"B1",x"38",x"30",x"06",x"20",x"58",x"B5",x"C8", -- 0x3538
    x"D0",x"F6",x"A4",x"3A",x"60",x"48",x"4A",x"4A", -- 0x3540
    x"4A",x"4A",x"20",x"50",x"B5",x"68",x"29",x"0F", -- 0x3548
    x"C9",x"0A",x"90",x"02",x"69",x"06",x"69",x"30", -- 0x3550
    x"C9",x"0D",x"D0",x"0B",x"20",x"EE",x"FF",x"4C", -- 0x3558
    x"28",x"BC",x"20",x"45",x"B5",x"A9",x"20",x"48", -- 0x3560
    x"A5",x"23",x"C5",x"1E",x"B0",x"03",x"20",x"25", -- 0x3568
    x"BC",x"68",x"E6",x"1E",x"6C",x"0E",x"02",x"25", -- 0x3570
    x"1F",x"F0",x"0E",x"8A",x"F0",x"0B",x"30",x"E5", -- 0x3578
    x"20",x"65",x"B5",x"20",x"58",x"B5",x"CA",x"D0", -- 0x3580
    x"F7",x"60",x"E6",x"0A",x"20",x"1D",x"9B",x"20", -- 0x3588
    x"4C",x"98",x"20",x"EE",x"92",x"A5",x"2A",x"85", -- 0x3590
    x"1F",x"4C",x"F6",x"8A",x"C8",x"B1",x"0B",x"C9", -- 0x3598
    x"4F",x"F0",x"E7",x"A9",x"00",x"85",x"3B",x"85", -- 0x35A0
    x"3C",x"20",x"D8",x"AE",x"20",x"DF",x"97",x"08", -- 0x35A8
    x"20",x"94",x"BD",x"A9",x"FF",x"85",x"2A",x"A9", -- 0x35B0
    x"7F",x"85",x"2B",x"28",x"90",x"11",x"20",x"97", -- 0x35B8
    x"8A",x"C9",x"2C",x"F0",x"13",x"20",x"EA",x"BD", -- 0x35C0
    x"20",x"94",x"BD",x"C6",x"0A",x"10",x"0C",x"20", -- 0x35C8
    x"97",x"8A",x"C9",x"2C",x"F0",x"02",x"C6",x"0A", -- 0x35D0
    x"20",x"DF",x"97",x"A5",x"2A",x"85",x"31",x"A5", -- 0x35D8
    x"2B",x"85",x"32",x"20",x"57",x"98",x"20",x"6F", -- 0x35E0
    x"BE",x"20",x"EA",x"BD",x"20",x"70",x"99",x"A5", -- 0x35E8
    x"3D",x"85",x"0B",x"A5",x"3E",x"85",x"0C",x"90", -- 0x35F0
    x"16",x"88",x"B0",x"06",x"20",x"25",x"BC",x"20", -- 0x35F8
    x"6D",x"98",x"B1",x"0B",x"85",x"2B",x"C8",x"B1", -- 0x3600
    x"0B",x"85",x"2A",x"C8",x"C8",x"84",x"0A",x"A5", -- 0x3608
    x"2A",x"18",x"E5",x"31",x"A5",x"2B",x"E5",x"32", -- 0x3610
    x"90",x"03",x"4C",x"F6",x"8A",x"20",x"23",x"99", -- 0x3618
    x"A2",x"FF",x"86",x"4D",x"A9",x"01",x"20",x"77", -- 0x3620
    x"B5",x"A6",x"3B",x"A9",x"02",x"20",x"77",x"B5", -- 0x3628
    x"A6",x"3C",x"A9",x"04",x"20",x"77",x"B5",x"A4", -- 0x3630
    x"0A",x"B1",x"0B",x"C9",x"0D",x"F0",x"BD",x"C9", -- 0x3638
    x"22",x"D0",x"0E",x"A9",x"FF",x"45",x"4D",x"85", -- 0x3640
    x"4D",x"A9",x"22",x"20",x"58",x"B5",x"C8",x"D0", -- 0x3648
    x"E8",x"24",x"4D",x"10",x"F6",x"C9",x"8D",x"D0", -- 0x3650
    x"0F",x"20",x"EB",x"97",x"84",x"0A",x"A9",x"00", -- 0x3658
    x"85",x"14",x"20",x"1F",x"99",x"4C",x"37",x"B6", -- 0x3660
    x"C9",x"E3",x"D0",x"02",x"E6",x"3B",x"C9",x"ED", -- 0x3668
    x"D0",x"06",x"A6",x"3B",x"F0",x"02",x"C6",x"3B", -- 0x3670
    x"C9",x"F5",x"D0",x"02",x"E6",x"3C",x"C9",x"FD", -- 0x3678
    x"D0",x"06",x"A6",x"3C",x"F0",x"02",x"C6",x"3C", -- 0x3680
    x"20",x"0E",x"B5",x"C8",x"D0",x"AB",x"00",x"20", -- 0x3688
    x"4E",x"6F",x"20",x"E3",x"00",x"20",x"C9",x"95", -- 0x3690
    x"D0",x"09",x"A6",x"26",x"F0",x"F0",x"B0",x"37", -- 0x3698
    x"4C",x"2A",x"98",x"B0",x"FB",x"A6",x"26",x"F0", -- 0x36A0
    x"E5",x"A5",x"2A",x"DD",x"F1",x"04",x"D0",x"0E", -- 0x36A8
    x"A5",x"2B",x"DD",x"F2",x"04",x"D0",x"07",x"A5", -- 0x36B0
    x"2C",x"DD",x"F3",x"04",x"F0",x"19",x"8A",x"38", -- 0x36B8
    x"E9",x"0F",x"AA",x"86",x"26",x"D0",x"E2",x"00", -- 0x36C0
    x"21",x"43",x"61",x"6E",x"27",x"74",x"20",x"4D", -- 0x36C8
    x"61",x"74",x"63",x"68",x"20",x"E3",x"00",x"BD", -- 0x36D0
    x"F1",x"04",x"85",x"2A",x"BD",x"F2",x"04",x"85", -- 0x36D8
    x"2B",x"BC",x"F3",x"04",x"C0",x"05",x"F0",x"7E", -- 0x36E0
    x"A0",x"00",x"B1",x"2A",x"7D",x"F4",x"04",x"91", -- 0x36E8
    x"2A",x"85",x"37",x"C8",x"B1",x"2A",x"7D",x"F5", -- 0x36F0
    x"04",x"91",x"2A",x"85",x"38",x"C8",x"B1",x"2A", -- 0x36F8
    x"7D",x"F6",x"04",x"91",x"2A",x"85",x"39",x"C8", -- 0x3700
    x"B1",x"2A",x"7D",x"F7",x"04",x"91",x"2A",x"A8", -- 0x3708
    x"A5",x"37",x"38",x"FD",x"F9",x"04",x"85",x"37", -- 0x3710
    x"A5",x"38",x"FD",x"FA",x"04",x"85",x"38",x"A5", -- 0x3718
    x"39",x"FD",x"FB",x"04",x"85",x"39",x"98",x"FD", -- 0x3720
    x"FC",x"04",x"05",x"37",x"05",x"38",x"05",x"39", -- 0x3728
    x"F0",x"0F",x"98",x"5D",x"F7",x"04",x"5D",x"FC", -- 0x3730
    x"04",x"10",x"04",x"B0",x"04",x"90",x"12",x"B0", -- 0x3738
    x"10",x"BC",x"FE",x"04",x"BD",x"FF",x"04",x"84", -- 0x3740
    x"0B",x"85",x"0C",x"20",x"77",x"98",x"4C",x"A3", -- 0x3748
    x"8B",x"A5",x"26",x"38",x"E9",x"0F",x"85",x"26", -- 0x3750
    x"A4",x"1B",x"84",x"0A",x"20",x"97",x"8A",x"C9", -- 0x3758
    x"2C",x"D0",x"3E",x"4C",x"95",x"B6",x"20",x"54", -- 0x3760
    x"B3",x"A5",x"26",x"18",x"69",x"F4",x"85",x"4B", -- 0x3768
    x"A9",x"05",x"85",x"4C",x"20",x"00",x"A5",x"A5", -- 0x3770
    x"2A",x"85",x"37",x"A5",x"2B",x"85",x"38",x"20", -- 0x3778
    x"E9",x"B4",x"A5",x"26",x"85",x"27",x"18",x"69", -- 0x3780
    x"F9",x"85",x"4B",x"A9",x"05",x"85",x"4C",x"20", -- 0x3788
    x"5F",x"9A",x"F0",x"AD",x"BD",x"F5",x"04",x"30", -- 0x3790
    x"04",x"B0",x"A6",x"90",x"B4",x"90",x"A2",x"B0", -- 0x3798
    x"B0",x"4C",x"96",x"8B",x"00",x"22",x"E3",x"20", -- 0x37A0
    x"76",x"61",x"72",x"69",x"61",x"62",x"6C",x"65", -- 0x37A8
    x"00",x"23",x"54",x"6F",x"6F",x"20",x"6D",x"61", -- 0x37B0
    x"6E",x"79",x"20",x"E3",x"73",x"00",x"24",x"4E", -- 0x37B8
    x"6F",x"20",x"B8",x"00",x"20",x"82",x"95",x"F0", -- 0x37C0
    x"DB",x"B0",x"D9",x"20",x"94",x"BD",x"20",x"41", -- 0x37C8
    x"98",x"20",x"B1",x"B4",x"A4",x"26",x"C0",x"96", -- 0x37D0
    x"B0",x"D6",x"A5",x"37",x"99",x"00",x"05",x"A5", -- 0x37D8
    x"38",x"99",x"01",x"05",x"A5",x"39",x"99",x"02", -- 0x37E0
    x"05",x"AA",x"20",x"8C",x"8A",x"C9",x"B8",x"D0", -- 0x37E8
    x"CC",x"E0",x"05",x"F0",x"5A",x"20",x"DD",x"92", -- 0x37F0
    x"A4",x"26",x"A5",x"2A",x"99",x"08",x"05",x"A5", -- 0x37F8
    x"2B",x"99",x"09",x"05",x"A5",x"2C",x"99",x"0A", -- 0x3800
    x"05",x"A5",x"2D",x"99",x"0B",x"05",x"A9",x"01", -- 0x3808
    x"20",x"D8",x"AE",x"20",x"8C",x"8A",x"C9",x"88", -- 0x3810
    x"D0",x"05",x"20",x"DD",x"92",x"A4",x"1B",x"84", -- 0x3818
    x"0A",x"A4",x"26",x"A5",x"2A",x"99",x"03",x"05", -- 0x3820
    x"A5",x"2B",x"99",x"04",x"05",x"A5",x"2C",x"99", -- 0x3828
    x"05",x"05",x"A5",x"2D",x"99",x"06",x"05",x"20", -- 0x3830
    x"80",x"98",x"A4",x"26",x"A5",x"0B",x"99",x"0D", -- 0x3838
    x"05",x"A5",x"0C",x"99",x"0E",x"05",x"18",x"98", -- 0x3840
    x"69",x"0F",x"85",x"26",x"4C",x"A3",x"8B",x"20", -- 0x3848
    x"29",x"9B",x"20",x"FD",x"92",x"A5",x"26",x"18", -- 0x3850
    x"69",x"08",x"85",x"4B",x"A9",x"05",x"85",x"4C", -- 0x3858
    x"20",x"8D",x"A3",x"20",x"99",x"A6",x"20",x"8C", -- 0x3860
    x"8A",x"C9",x"88",x"D0",x"08",x"20",x"29",x"9B", -- 0x3868
    x"20",x"FD",x"92",x"A4",x"1B",x"84",x"0A",x"A5", -- 0x3870
    x"26",x"18",x"69",x"03",x"85",x"4B",x"A9",x"05", -- 0x3878
    x"85",x"4C",x"20",x"8D",x"A3",x"4C",x"37",x"B8", -- 0x3880
    x"20",x"9A",x"B9",x"20",x"57",x"98",x"A4",x"25", -- 0x3888
    x"C0",x"1A",x"B0",x"0E",x"A5",x"0B",x"99",x"CC", -- 0x3890
    x"05",x"A5",x"0C",x"99",x"E6",x"05",x"E6",x"25", -- 0x3898
    x"90",x"30",x"00",x"25",x"54",x"6F",x"6F",x"20", -- 0x38A0
    x"6D",x"61",x"6E",x"79",x"20",x"E4",x"73",x"00", -- 0x38A8
    x"26",x"4E",x"6F",x"20",x"E4",x"00",x"20",x"57", -- 0x38B0
    x"98",x"A6",x"25",x"F0",x"F2",x"C6",x"25",x"BC", -- 0x38B8
    x"CB",x"05",x"BD",x"E5",x"05",x"84",x"0B",x"85", -- 0x38C0
    x"0C",x"4C",x"9B",x"8B",x"20",x"9A",x"B9",x"20", -- 0x38C8
    x"57",x"98",x"A5",x"20",x"F0",x"03",x"20",x"05", -- 0x38D0
    x"99",x"A4",x"3D",x"A5",x"3E",x"84",x"0B",x"85", -- 0x38D8
    x"0C",x"4C",x"A3",x"8B",x"20",x"57",x"98",x"A9", -- 0x38E0
    x"33",x"85",x"16",x"A9",x"B4",x"85",x"17",x"4C", -- 0x38E8
    x"9B",x"8B",x"20",x"97",x"8A",x"C9",x"87",x"F0", -- 0x38F0
    x"EB",x"A4",x"0A",x"88",x"20",x"6D",x"98",x"A5", -- 0x38F8
    x"0B",x"85",x"16",x"A5",x"0C",x"85",x"17",x"4C", -- 0x3900
    x"7D",x"8B",x"00",x"27",x"EE",x"20",x"73",x"79", -- 0x3908
    x"6E",x"74",x"61",x"78",x"00",x"20",x"97",x"8A", -- 0x3910
    x"C9",x"85",x"F0",x"D6",x"C6",x"0A",x"20",x"1D", -- 0x3918
    x"9B",x"20",x"F0",x"92",x"A4",x"1B",x"C8",x"84", -- 0x3920
    x"0A",x"E0",x"E5",x"F0",x"04",x"E0",x"E4",x"D0", -- 0x3928
    x"D9",x"8A",x"48",x"A5",x"2B",x"05",x"2C",x"05", -- 0x3930
    x"2D",x"D0",x"42",x"A6",x"2A",x"F0",x"3E",x"CA", -- 0x3938
    x"F0",x"1A",x"A4",x"0A",x"B1",x"0B",x"C8",x"C9", -- 0x3940
    x"0D",x"F0",x"32",x"C9",x"3A",x"F0",x"2E",x"C9", -- 0x3948
    x"8B",x"F0",x"2A",x"C9",x"2C",x"D0",x"ED",x"CA", -- 0x3950
    x"D0",x"EA",x"84",x"0A",x"20",x"9A",x"B9",x"68", -- 0x3958
    x"C9",x"E4",x"F0",x"06",x"20",x"77",x"98",x"4C", -- 0x3960
    x"D2",x"B8",x"A4",x"0A",x"B1",x"0B",x"C8",x"C9", -- 0x3968
    x"0D",x"F0",x"04",x"C9",x"3A",x"D0",x"F5",x"88", -- 0x3970
    x"84",x"0A",x"4C",x"8B",x"B8",x"A4",x"0A",x"68", -- 0x3978
    x"B1",x"0B",x"C8",x"C9",x"8B",x"F0",x"0E",x"C9", -- 0x3980
    x"0D",x"D0",x"F5",x"00",x"28",x"EE",x"20",x"72", -- 0x3988
    x"61",x"6E",x"67",x"65",x"00",x"84",x"0A",x"4C", -- 0x3990
    x"E3",x"98",x"20",x"DF",x"97",x"B0",x"10",x"20", -- 0x3998
    x"1D",x"9B",x"20",x"F0",x"92",x"A5",x"1B",x"85", -- 0x39A0
    x"0A",x"A5",x"2B",x"29",x"7F",x"85",x"2B",x"20", -- 0x39A8
    x"70",x"99",x"B0",x"01",x"60",x"00",x"29",x"4E", -- 0x39B0
    x"6F",x"20",x"73",x"75",x"63",x"68",x"20",x"6C", -- 0x39B8
    x"69",x"6E",x"65",x"00",x"4C",x"0E",x"8C",x"4C", -- 0x39C0
    x"2A",x"98",x"84",x"0A",x"4C",x"98",x"8B",x"C6", -- 0x39C8
    x"0A",x"20",x"A9",x"BF",x"A5",x"1B",x"85",x"0A", -- 0x39D0
    x"84",x"4D",x"20",x"97",x"8A",x"C9",x"2C",x"D0", -- 0x39D8
    x"E9",x"A5",x"4D",x"48",x"20",x"82",x"95",x"F0", -- 0x39E0
    x"DE",x"A5",x"1B",x"85",x"0A",x"68",x"85",x"4D", -- 0x39E8
    x"08",x"20",x"94",x"BD",x"A4",x"4D",x"20",x"D7", -- 0x39F0
    x"FF",x"85",x"27",x"28",x"90",x"1B",x"A5",x"27", -- 0x39F8
    x"D0",x"C2",x"20",x"D7",x"FF",x"85",x"36",x"AA", -- 0x3A00
    x"F0",x"09",x"20",x"D7",x"FF",x"9D",x"FF",x"05", -- 0x3A08
    x"CA",x"D0",x"F7",x"20",x"1E",x"8C",x"4C",x"DA", -- 0x3A10
    x"B9",x"A5",x"27",x"F0",x"A7",x"30",x"0C",x"A2", -- 0x3A18
    x"03",x"20",x"D7",x"FF",x"95",x"2A",x"CA",x"10", -- 0x3A20
    x"F8",x"30",x"0E",x"A2",x"04",x"20",x"D7",x"FF", -- 0x3A28
    x"9D",x"6C",x"04",x"CA",x"10",x"F7",x"20",x"B2", -- 0x3A30
    x"A3",x"20",x"B4",x"B4",x"4C",x"DA",x"B9",x"68", -- 0x3A38
    x"68",x"4C",x"98",x"8B",x"20",x"97",x"8A",x"C9", -- 0x3A40
    x"23",x"F0",x"84",x"C9",x"86",x"F0",x"03",x"C6", -- 0x3A48
    x"0A",x"18",x"66",x"4D",x"46",x"4D",x"A9",x"FF", -- 0x3A50
    x"85",x"4E",x"20",x"8A",x"8E",x"B0",x"0A",x"20", -- 0x3A58
    x"8A",x"8E",x"90",x"FB",x"A2",x"FF",x"86",x"4E", -- 0x3A60
    x"18",x"08",x"06",x"4D",x"28",x"66",x"4D",x"C9", -- 0x3A68
    x"2C",x"F0",x"E7",x"C9",x"3B",x"F0",x"E3",x"C6", -- 0x3A70
    x"0A",x"A5",x"4D",x"48",x"A5",x"4E",x"48",x"20", -- 0x3A78
    x"82",x"95",x"F0",x"BB",x"68",x"85",x"4E",x"68", -- 0x3A80
    x"85",x"4D",x"A5",x"1B",x"85",x"0A",x"08",x"24", -- 0x3A88
    x"4D",x"70",x"06",x"A5",x"4E",x"C9",x"FF",x"D0", -- 0x3A90
    x"17",x"24",x"4D",x"10",x"05",x"A9",x"3F",x"20", -- 0x3A98
    x"58",x"B5",x"20",x"FC",x"BB",x"84",x"36",x"06", -- 0x3AA0
    x"4D",x"18",x"66",x"4D",x"24",x"4D",x"70",x"1D", -- 0x3AA8
    x"85",x"1B",x"A9",x"00",x"85",x"19",x"A9",x"06", -- 0x3AB0
    x"85",x"1A",x"20",x"AD",x"AD",x"20",x"8C",x"8A", -- 0x3AB8
    x"C9",x"2C",x"F0",x"06",x"C9",x"0D",x"D0",x"F5", -- 0x3AC0
    x"A0",x"FE",x"C8",x"84",x"4E",x"28",x"B0",x"0C", -- 0x3AC8
    x"20",x"94",x"BD",x"20",x"34",x"AC",x"20",x"B4", -- 0x3AD0
    x"B4",x"4C",x"5A",x"BA",x"A9",x"00",x"85",x"27", -- 0x3AD8
    x"20",x"21",x"8C",x"4C",x"5A",x"BA",x"A0",x"00", -- 0x3AE0
    x"84",x"3D",x"A4",x"18",x"84",x"3E",x"20",x"97", -- 0x3AE8
    x"8A",x"C6",x"0A",x"C9",x"3A",x"F0",x"10",x"C9", -- 0x3AF0
    x"0D",x"F0",x"0C",x"C9",x"8B",x"F0",x"08",x"20", -- 0x3AF8
    x"9A",x"B9",x"A0",x"01",x"20",x"55",x"BE",x"20", -- 0x3B00
    x"57",x"98",x"A5",x"3D",x"85",x"1C",x"A5",x"3E", -- 0x3B08
    x"85",x"1D",x"4C",x"9B",x"8B",x"20",x"97",x"8A", -- 0x3B10
    x"C9",x"2C",x"F0",x"03",x"4C",x"96",x"8B",x"20", -- 0x3B18
    x"82",x"95",x"F0",x"F1",x"B0",x"0C",x"20",x"50", -- 0x3B20
    x"BB",x"20",x"94",x"BD",x"20",x"B1",x"B4",x"4C", -- 0x3B28
    x"40",x"BB",x"20",x"50",x"BB",x"20",x"94",x"BD", -- 0x3B30
    x"20",x"AD",x"AD",x"85",x"27",x"20",x"1E",x"8C", -- 0x3B38
    x"18",x"A5",x"1B",x"65",x"19",x"85",x"1C",x"A5", -- 0x3B40
    x"1A",x"69",x"00",x"85",x"1D",x"4C",x"15",x"BB", -- 0x3B48
    x"A5",x"1B",x"85",x"0A",x"A5",x"1C",x"85",x"19", -- 0x3B50
    x"A5",x"1D",x"85",x"1A",x"A0",x"00",x"84",x"1B", -- 0x3B58
    x"20",x"8C",x"8A",x"C9",x"2C",x"F0",x"49",x"C9", -- 0x3B60
    x"DC",x"F0",x"45",x"C9",x"0D",x"F0",x"0B",x"20", -- 0x3B68
    x"8C",x"8A",x"C9",x"2C",x"F0",x"3A",x"C9",x"0D", -- 0x3B70
    x"D0",x"F5",x"A4",x"1B",x"B1",x"19",x"30",x"1C", -- 0x3B78
    x"C8",x"C8",x"B1",x"19",x"AA",x"C8",x"B1",x"19", -- 0x3B80
    x"C9",x"20",x"F0",x"F9",x"C9",x"DC",x"F0",x"1D", -- 0x3B88
    x"8A",x"18",x"65",x"19",x"85",x"19",x"90",x"E2", -- 0x3B90
    x"E6",x"1A",x"B0",x"DE",x"00",x"2A",x"4F",x"75", -- 0x3B98
    x"74",x"20",x"6F",x"66",x"20",x"DC",x"00",x"2B", -- 0x3BA0
    x"4E",x"6F",x"20",x"F5",x"00",x"C8",x"84",x"1B", -- 0x3BA8
    x"60",x"20",x"1D",x"9B",x"20",x"4C",x"98",x"20", -- 0x3BB0
    x"EE",x"92",x"A6",x"24",x"F0",x"E8",x"A5",x"2A", -- 0x3BB8
    x"05",x"2B",x"05",x"2C",x"05",x"2D",x"F0",x"05", -- 0x3BC0
    x"C6",x"24",x"4C",x"9B",x"8B",x"BC",x"A3",x"05", -- 0x3BC8
    x"BD",x"B7",x"05",x"4C",x"DD",x"B8",x"00",x"2C", -- 0x3BD0
    x"54",x"6F",x"6F",x"20",x"6D",x"61",x"6E",x"79", -- 0x3BD8
    x"20",x"F5",x"73",x"00",x"A6",x"24",x"E0",x"14", -- 0x3BE0
    x"B0",x"EC",x"20",x"6D",x"98",x"A5",x"0B",x"9D", -- 0x3BE8
    x"A4",x"05",x"A5",x"0C",x"9D",x"B8",x"05",x"E6", -- 0x3BF0
    x"24",x"4C",x"A3",x"8B",x"A0",x"00",x"A9",x"06", -- 0x3BF8
    x"D0",x"07",x"20",x"58",x"B5",x"A0",x"00",x"A9", -- 0x3C00
    x"07",x"84",x"37",x"85",x"38",x"A9",x"EE",x"85", -- 0x3C08
    x"39",x"A9",x"20",x"85",x"3A",x"A0",x"FF",x"84", -- 0x3C10
    x"3B",x"C8",x"A2",x"37",x"98",x"20",x"F1",x"FF", -- 0x3C18
    x"90",x"06",x"4C",x"38",x"98",x"20",x"E7",x"FF", -- 0x3C20
    x"A9",x"00",x"85",x"1E",x"60",x"20",x"70",x"99", -- 0x3C28
    x"B0",x"4E",x"A5",x"3D",x"E9",x"02",x"85",x"37", -- 0x3C30
    x"85",x"3D",x"85",x"12",x"A5",x"3E",x"E9",x"00", -- 0x3C38
    x"85",x"38",x"85",x"13",x"85",x"3E",x"A0",x"03", -- 0x3C40
    x"B1",x"37",x"18",x"65",x"37",x"85",x"37",x"90", -- 0x3C48
    x"02",x"E6",x"38",x"A0",x"00",x"B1",x"37",x"91", -- 0x3C50
    x"12",x"C9",x"0D",x"F0",x"09",x"C8",x"D0",x"F5", -- 0x3C58
    x"E6",x"38",x"E6",x"13",x"D0",x"EF",x"C8",x"D0", -- 0x3C60
    x"04",x"E6",x"38",x"E6",x"13",x"B1",x"37",x"91", -- 0x3C68
    x"12",x"30",x"09",x"20",x"81",x"BC",x"20",x"81", -- 0x3C70
    x"BC",x"4C",x"5D",x"BC",x"20",x"92",x"BE",x"18", -- 0x3C78
    x"60",x"C8",x"D0",x"04",x"E6",x"13",x"E6",x"38", -- 0x3C80
    x"B1",x"37",x"91",x"12",x"60",x"84",x"3B",x"20", -- 0x3C88
    x"2D",x"BC",x"A0",x"07",x"84",x"3C",x"A0",x"00", -- 0x3C90
    x"A9",x"0D",x"D1",x"3B",x"F0",x"72",x"C8",x"D1", -- 0x3C98
    x"3B",x"D0",x"FB",x"C8",x"C8",x"C8",x"84",x"3F", -- 0x3CA0
    x"E6",x"3F",x"A5",x"12",x"85",x"39",x"A5",x"13", -- 0x3CA8
    x"85",x"3A",x"20",x"92",x"BE",x"85",x"37",x"A5", -- 0x3CB0
    x"13",x"85",x"38",x"88",x"A5",x"06",x"C5",x"12", -- 0x3CB8
    x"A5",x"07",x"E5",x"13",x"B0",x"10",x"20",x"6F", -- 0x3CC0
    x"BE",x"20",x"20",x"BD",x"00",x"00",x"86",x"20", -- 0x3CC8
    x"73",x"70",x"61",x"63",x"65",x"00",x"B1",x"39", -- 0x3CD0
    x"91",x"37",x"98",x"D0",x"04",x"C6",x"3A",x"C6", -- 0x3CD8
    x"38",x"88",x"98",x"65",x"39",x"A6",x"3A",x"90", -- 0x3CE0
    x"01",x"E8",x"C5",x"3D",x"8A",x"E5",x"3E",x"B0", -- 0x3CE8
    x"E5",x"38",x"A0",x"01",x"A5",x"2B",x"91",x"3D", -- 0x3CF0
    x"C8",x"A5",x"2A",x"91",x"3D",x"C8",x"A5",x"3F", -- 0x3CF8
    x"91",x"3D",x"20",x"56",x"BE",x"A0",x"FF",x"C8", -- 0x3D00
    x"B1",x"3B",x"91",x"3D",x"C9",x"0D",x"D0",x"F7", -- 0x3D08
    x"60",x"20",x"57",x"98",x"20",x"20",x"BD",x"A5", -- 0x3D10
    x"18",x"85",x"0C",x"86",x"0B",x"4C",x"0B",x"8B", -- 0x3D18
    x"A5",x"12",x"85",x"00",x"85",x"02",x"A5",x"13", -- 0x3D20
    x"85",x"01",x"85",x"03",x"20",x"3A",x"BD",x"A2", -- 0x3D28
    x"80",x"A9",x"00",x"9D",x"7F",x"04",x"CA",x"D0", -- 0x3D30
    x"FA",x"60",x"A5",x"18",x"85",x"1D",x"A5",x"06", -- 0x3D38
    x"85",x"04",x"A5",x"07",x"85",x"05",x"A9",x"00", -- 0x3D40
    x"85",x"24",x"85",x"26",x"85",x"25",x"85",x"1C", -- 0x3D48
    x"60",x"A5",x"04",x"38",x"E9",x"05",x"20",x"2E", -- 0x3D50
    x"BE",x"A0",x"00",x"A5",x"30",x"91",x"04",x"C8", -- 0x3D58
    x"A5",x"2E",x"29",x"80",x"85",x"2E",x"A5",x"31", -- 0x3D60
    x"29",x"7F",x"05",x"2E",x"91",x"04",x"C8",x"A5", -- 0x3D68
    x"32",x"91",x"04",x"C8",x"A5",x"33",x"91",x"04", -- 0x3D70
    x"C8",x"A5",x"34",x"91",x"04",x"60",x"A5",x"04", -- 0x3D78
    x"18",x"85",x"4B",x"69",x"05",x"85",x"04",x"A5", -- 0x3D80
    x"05",x"85",x"4C",x"69",x"00",x"85",x"05",x"60", -- 0x3D88
    x"F0",x"20",x"30",x"BD",x"A5",x"04",x"38",x"E9", -- 0x3D90
    x"04",x"20",x"2E",x"BE",x"A0",x"03",x"A5",x"2D", -- 0x3D98
    x"91",x"04",x"88",x"A5",x"2C",x"91",x"04",x"88", -- 0x3DA0
    x"A5",x"2B",x"91",x"04",x"88",x"A5",x"2A",x"91", -- 0x3DA8
    x"04",x"60",x"18",x"A5",x"04",x"E5",x"36",x"20", -- 0x3DB0
    x"2E",x"BE",x"A4",x"36",x"F0",x"08",x"B9",x"FF", -- 0x3DB8
    x"05",x"91",x"04",x"88",x"D0",x"F8",x"A5",x"36", -- 0x3DC0
    x"91",x"04",x"60",x"A0",x"00",x"B1",x"04",x"85", -- 0x3DC8
    x"36",x"F0",x"09",x"A8",x"B1",x"04",x"99",x"FF", -- 0x3DD0
    x"05",x"88",x"D0",x"F8",x"A0",x"00",x"B1",x"04", -- 0x3DD8
    x"38",x"65",x"04",x"85",x"04",x"90",x"23",x"E6", -- 0x3DE0
    x"05",x"60",x"A0",x"03",x"B1",x"04",x"85",x"2D", -- 0x3DE8
    x"88",x"B1",x"04",x"85",x"2C",x"88",x"B1",x"04", -- 0x3DF0
    x"85",x"2B",x"88",x"B1",x"04",x"85",x"2A",x"18", -- 0x3DF8
    x"A5",x"04",x"69",x"04",x"85",x"04",x"90",x"02", -- 0x3E00
    x"E6",x"05",x"60",x"A2",x"37",x"A0",x"03",x"B1", -- 0x3E08
    x"04",x"95",x"03",x"88",x"B1",x"04",x"95",x"02", -- 0x3E10
    x"88",x"B1",x"04",x"95",x"01",x"88",x"B1",x"04", -- 0x3E18
    x"95",x"00",x"18",x"A5",x"04",x"69",x"04",x"85", -- 0x3E20
    x"04",x"90",x"DF",x"E6",x"05",x"60",x"85",x"04", -- 0x3E28
    x"B0",x"02",x"C6",x"05",x"A4",x"05",x"C4",x"03", -- 0x3E30
    x"90",x"07",x"D0",x"04",x"C5",x"02",x"90",x"01", -- 0x3E38
    x"60",x"4C",x"B7",x"8C",x"A5",x"2A",x"95",x"00", -- 0x3E40
    x"A5",x"2B",x"95",x"01",x"A5",x"2C",x"95",x"02", -- 0x3E48
    x"A5",x"2D",x"95",x"03",x"60",x"18",x"98",x"65", -- 0x3E50
    x"3D",x"85",x"3D",x"90",x"02",x"E6",x"3E",x"A0", -- 0x3E58
    x"01",x"60",x"20",x"DD",x"BE",x"A8",x"A9",x"FF", -- 0x3E60
    x"84",x"3D",x"A2",x"37",x"20",x"DD",x"FF",x"A5", -- 0x3E68
    x"18",x"85",x"13",x"A0",x"00",x"84",x"12",x"C8", -- 0x3E70
    x"88",x"B1",x"12",x"C9",x"0D",x"D0",x"1F",x"C8", -- 0x3E78
    x"B1",x"12",x"30",x"0C",x"A0",x"03",x"B1",x"12", -- 0x3E80
    x"F0",x"14",x"18",x"20",x"93",x"BE",x"D0",x"E8", -- 0x3E88
    x"C8",x"18",x"98",x"65",x"12",x"85",x"12",x"90", -- 0x3E90
    x"02",x"E6",x"13",x"A0",x"01",x"60",x"20",x"CF", -- 0x3E98
    x"BF",x"0D",x"42",x"61",x"64",x"20",x"70",x"72", -- 0x3EA0
    x"6F",x"67",x"72",x"61",x"6D",x"0D",x"EA",x"4C", -- 0x3EA8
    x"F6",x"8A",x"A9",x"00",x"85",x"37",x"A9",x"06", -- 0x3EB0
    x"85",x"38",x"A4",x"36",x"A9",x"0D",x"99",x"00", -- 0x3EB8
    x"06",x"60",x"20",x"D2",x"BE",x"A2",x"00",x"A0", -- 0x3EC0
    x"06",x"20",x"F7",x"FF",x"4C",x"9B",x"8B",x"4C", -- 0x3EC8
    x"0E",x"8C",x"20",x"1D",x"9B",x"D0",x"F8",x"20", -- 0x3ED0
    x"B2",x"BE",x"4C",x"4C",x"98",x"20",x"D2",x"BE", -- 0x3ED8
    x"88",x"84",x"39",x"A5",x"18",x"85",x"3A",x"A9", -- 0x3EE0
    x"82",x"20",x"F4",x"FF",x"86",x"3B",x"84",x"3C", -- 0x3EE8
    x"A9",x"00",x"60",x"20",x"6F",x"BE",x"A5",x"12", -- 0x3EF0
    x"85",x"45",x"A5",x"13",x"85",x"46",x"A9",x"23", -- 0x3EF8
    x"85",x"3D",x"A9",x"80",x"85",x"3E",x"A5",x"18", -- 0x3F00
    x"85",x"42",x"20",x"DD",x"BE",x"86",x"3F",x"84", -- 0x3F08
    x"40",x"86",x"43",x"84",x"44",x"86",x"47",x"84", -- 0x3F10
    x"48",x"85",x"41",x"A8",x"A2",x"37",x"20",x"DD", -- 0x3F18
    x"FF",x"4C",x"9B",x"8B",x"20",x"62",x"BE",x"4C", -- 0x3F20
    x"F3",x"8A",x"20",x"62",x"BE",x"4C",x"14",x"BD", -- 0x3F28
    x"20",x"A9",x"BF",x"48",x"20",x"13",x"98",x"20", -- 0x3F30
    x"EE",x"92",x"68",x"A8",x"A2",x"2A",x"A9",x"01", -- 0x3F38
    x"20",x"DA",x"FF",x"4C",x"9B",x"8B",x"38",x"A9", -- 0x3F40
    x"00",x"2A",x"2A",x"48",x"20",x"B5",x"BF",x"A2", -- 0x3F48
    x"2A",x"68",x"20",x"DA",x"FF",x"A9",x"40",x"60", -- 0x3F50
    x"20",x"A9",x"BF",x"48",x"20",x"AE",x"8A",x"20", -- 0x3F58
    x"49",x"98",x"20",x"EE",x"92",x"68",x"A8",x"A5", -- 0x3F60
    x"2A",x"20",x"D4",x"FF",x"4C",x"9B",x"8B",x"20", -- 0x3F68
    x"B5",x"BF",x"20",x"D7",x"FF",x"4C",x"D8",x"AE", -- 0x3F70
    x"A9",x"40",x"D0",x"06",x"A9",x"80",x"D0",x"02", -- 0x3F78
    x"A9",x"C0",x"48",x"20",x"EC",x"AD",x"D0",x"0E", -- 0x3F80
    x"20",x"BA",x"BE",x"A2",x"00",x"A0",x"06",x"68", -- 0x3F88
    x"20",x"CE",x"FF",x"4C",x"D8",x"AE",x"4C",x"0E", -- 0x3F90
    x"8C",x"20",x"A9",x"BF",x"20",x"52",x"98",x"A4", -- 0x3F98
    x"2A",x"A9",x"00",x"20",x"CE",x"FF",x"4C",x"9B", -- 0x3FA0
    x"8B",x"A5",x"0A",x"85",x"1B",x"A5",x"0B",x"85", -- 0x3FA8
    x"19",x"A5",x"0C",x"85",x"1A",x"20",x"8C",x"8A", -- 0x3FB0
    x"C9",x"23",x"D0",x"07",x"20",x"E3",x"92",x"A4", -- 0x3FB8
    x"2A",x"98",x"60",x"00",x"2D",x"4D",x"69",x"73", -- 0x3FC0
    x"73",x"69",x"6E",x"67",x"20",x"23",x"00",x"68", -- 0x3FC8
    x"85",x"37",x"68",x"85",x"38",x"A0",x"00",x"F0", -- 0x3FD0
    x"03",x"20",x"E3",x"FF",x"20",x"4B",x"89",x"10", -- 0x3FD8
    x"F8",x"6C",x"37",x"00",x"20",x"57",x"98",x"20", -- 0x3FE0
    x"25",x"BC",x"A0",x"01",x"B1",x"FD",x"F0",x"06", -- 0x3FE8
    x"20",x"0E",x"B5",x"C8",x"D0",x"F6",x"4C",x"9B", -- 0x3FF0
    x"8B",x"00",x"52",x"6F",x"67",x"65",x"72",x"00"  -- 0x3FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
     DATA <= ROM(to_integer(unsigned(ADDR)));
  end process;
end RTL;
