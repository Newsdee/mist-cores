-- generated with romgen by MikeJ
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity BBC_SUPERMMC_ROM is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of BBC_SUPERMMC_ROM is


  type ROM_ARRAY is array(0 to 16383) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"00",x"00",x"00",x"4C",x"55",x"94",x"82",x"11", -- 0x0000
    x"5A",x"44",x"46",x"53",x"00",x"30",x"2E",x"39", -- 0x0008
    x"30",x"00",x"28",x"43",x"29",x"6C",x"1E",x"02", -- 0x0010
    x"20",x"5B",x"80",x"44",x"69",x"73",x"6B",x"20", -- 0x0018
    x"90",x"11",x"20",x"5B",x"80",x"42",x"61",x"64", -- 0x0020
    x"20",x"90",x"08",x"20",x"5B",x"80",x"46",x"69", -- 0x0028
    x"6C",x"65",x"20",x"85",x"B3",x"68",x"85",x"AE", -- 0x0030
    x"68",x"85",x"AF",x"A5",x"B3",x"48",x"98",x"48", -- 0x0038
    x"A0",x"00",x"20",x"DA",x"83",x"B1",x"AE",x"8D", -- 0x0040
    x"01",x"01",x"2C",x"DE",x"10",x"10",x"25",x"A9", -- 0x0048
    x"02",x"8D",x"DE",x"10",x"A9",x"00",x"8D",x"00", -- 0x0050
    x"01",x"F0",x"19",x"A9",x"02",x"8D",x"DE",x"10", -- 0x0058
    x"A9",x"00",x"8D",x"00",x"01",x"85",x"B3",x"68", -- 0x0060
    x"85",x"AE",x"68",x"85",x"AF",x"A5",x"B3",x"48", -- 0x0068
    x"98",x"48",x"A0",x"00",x"20",x"DA",x"83",x"B1", -- 0x0070
    x"AE",x"30",x"08",x"F0",x"0D",x"20",x"9C",x"80", -- 0x0078
    x"4C",x"74",x"80",x"68",x"A8",x"68",x"18",x"6C", -- 0x0080
    x"AE",x"00",x"A9",x"00",x"AE",x"DE",x"10",x"9D", -- 0x0088
    x"00",x"01",x"A9",x"FF",x"8D",x"DE",x"10",x"4C", -- 0x0090
    x"00",x"01",x"A9",x"2E",x"20",x"E1",x"83",x"2C", -- 0x0098
    x"DE",x"10",x"10",x"14",x"48",x"20",x"1C",x"99", -- 0x00A0
    x"8A",x"48",x"09",x"10",x"20",x"17",x"99",x"68", -- 0x00A8
    x"AA",x"68",x"20",x"E3",x"FF",x"4C",x"18",x"99", -- 0x00B0
    x"AE",x"DE",x"10",x"9D",x"00",x"01",x"EE",x"DE", -- 0x00B8
    x"10",x"60",x"48",x"20",x"05",x"82",x"20",x"CA", -- 0x00C0
    x"80",x"68",x"48",x"29",x"0F",x"C9",x"0A",x"90", -- 0x00C8
    x"02",x"69",x"06",x"69",x"30",x"20",x"9C",x"80", -- 0x00D0
    x"68",x"60",x"20",x"EA",x"80",x"CA",x"CA",x"20", -- 0x00D8
    x"E2",x"80",x"B1",x"B0",x"9D",x"72",x"10",x"E8", -- 0x00E0
    x"C8",x"60",x"20",x"ED",x"80",x"B1",x"B0",x"95", -- 0x00E8
    x"BC",x"E8",x"C8",x"60",x"A9",x"20",x"A2",x"06", -- 0x00F0
    x"95",x"C7",x"CA",x"10",x"FB",x"60",x"20",x"4D", -- 0x00F8
    x"83",x"20",x"F4",x"80",x"30",x"13",x"20",x"4D", -- 0x0100
    x"83",x"20",x"F4",x"80",x"A5",x"BC",x"85",x"F2", -- 0x0108
    x"A5",x"BD",x"85",x"F3",x"A0",x"00",x"20",x"BF", -- 0x0110
    x"86",x"A2",x"01",x"20",x"C5",x"FF",x"B0",x"DD", -- 0x0118
    x"85",x"C7",x"C9",x"2E",x"D0",x"04",x"A9",x"20", -- 0x0120
    x"D0",x"4D",x"C9",x"3A",x"D0",x"21",x"20",x"C5", -- 0x0128
    x"FF",x"B0",x"15",x"38",x"E9",x"30",x"90",x"10", -- 0x0130
    x"C9",x"04",x"B0",x"0C",x"20",x"7E",x"87",x"20", -- 0x0138
    x"C5",x"FF",x"B0",x"5C",x"C9",x"2E",x"F0",x"03", -- 0x0140
    x"4C",x"74",x"83",x"A9",x"24",x"D0",x"28",x"C9", -- 0x0148
    x"2A",x"D0",x"19",x"20",x"C5",x"FF",x"B0",x"08", -- 0x0150
    x"C9",x"2E",x"D0",x"32",x"A9",x"23",x"D0",x"17", -- 0x0158
    x"A2",x"00",x"A9",x"23",x"95",x"C7",x"E8",x"E0", -- 0x0160
    x"07",x"D0",x"F9",x"60",x"20",x"C5",x"FF",x"B0", -- 0x0168
    x"2F",x"C9",x"2E",x"D0",x"10",x"A5",x"C7",x"85", -- 0x0170
    x"CE",x"4C",x"1B",x"81",x"20",x"C5",x"FF",x"B0", -- 0x0178
    x"1F",x"E0",x"07",x"F0",x"09",x"C9",x"2A",x"D0", -- 0x0180
    x"12",x"20",x"C5",x"FF",x"B0",x"D4",x"20",x"22", -- 0x0188
    x"80",x"CC",x"66",x"69",x"6C",x"65",x"6E",x"61", -- 0x0190
    x"6D",x"65",x"00",x"95",x"C7",x"E8",x"D0",x"DC", -- 0x0198
    x"60",x"20",x"E1",x"83",x"AD",x"04",x"0F",x"20", -- 0x01A0
    x"47",x"83",x"CD",x"04",x"0F",x"F0",x"F1",x"20", -- 0x01A8
    x"33",x"80",x"C8",x"44",x"69",x"73",x"6B",x"20", -- 0x01B0
    x"63",x"68",x"61",x"6E",x"67",x"65",x"64",x"00", -- 0x01B8
    x"20",x"E1",x"83",x"B9",x"0F",x"0E",x"08",x"29", -- 0x01C0
    x"7F",x"D0",x"05",x"20",x"CB",x"9F",x"F0",x"06", -- 0x01C8
    x"20",x"9C",x"80",x"20",x"9A",x"80",x"A2",x"06", -- 0x01D0
    x"B9",x"08",x"0E",x"29",x"7F",x"20",x"9C",x"80", -- 0x01D8
    x"C8",x"CA",x"10",x"F4",x"20",x"CB",x"9F",x"A9", -- 0x01E0
    x"20",x"28",x"10",x"02",x"A9",x"4C",x"20",x"9C", -- 0x01E8
    x"80",x"4C",x"CE",x"9F",x"20",x"CE",x"9F",x"88", -- 0x01F0
    x"D0",x"FA",x"60",x"4A",x"4A",x"4A",x"4A",x"4A", -- 0x01F8
    x"4A",x"29",x"03",x"60",x"4A",x"4A",x"4A",x"4A", -- 0x0200
    x"4A",x"60",x"0A",x"0A",x"0A",x"0A",x"0A",x"60", -- 0x0208
    x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8", -- 0x0210
    x"60",x"88",x"88",x"88",x"88",x"88",x"88",x"88", -- 0x0218
    x"88",x"60",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0220
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0228
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0230
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0238
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0240
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0248
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0250
    x"00",x"00",x"00",x"00",x"00",x"60",x"A9",x"23", -- 0x0258
    x"D0",x"02",x"A9",x"FF",x"8D",x"CF",x"10",x"60", -- 0x0260
    x"20",x"FE",x"80",x"4C",x"71",x"82",x"20",x"06", -- 0x0268
    x"81",x"20",x"96",x"82",x"B0",x"E7",x"20",x"2B", -- 0x0270
    x"80",x"D6",x"6E",x"6F",x"74",x"20",x"66",x"6F", -- 0x0278
    x"75",x"6E",x"64",x"00",x"20",x"5E",x"82",x"20", -- 0x0280
    x"01",x"9A",x"20",x"68",x"82",x"20",x"01",x"83", -- 0x0288
    x"20",x"9D",x"82",x"B0",x"F8",x"60",x"20",x"4D", -- 0x0290
    x"AB",x"A0",x"F8",x"D0",x"03",x"AC",x"CE",x"10", -- 0x0298
    x"20",x"10",x"82",x"CC",x"05",x"0F",x"B0",x"44", -- 0x02A0
    x"20",x"10",x"82",x"A2",x"07",x"B5",x"C7",x"CD", -- 0x02A8
    x"CF",x"10",x"F0",x"0E",x"20",x"EE",x"82",x"59", -- 0x02B0
    x"07",x"0E",x"B0",x"02",x"29",x"DF",x"29",x"7F", -- 0x02B8
    x"D0",x"09",x"88",x"CA",x"10",x"E7",x"8C",x"CE", -- 0x02C0
    x"10",x"38",x"60",x"88",x"CA",x"10",x"FC",x"30", -- 0x02C8
    x"CF",x"20",x"4C",x"98",x"B9",x"10",x"0E",x"99", -- 0x02D0
    x"08",x"0E",x"B9",x"10",x"0F",x"99",x"08",x"0F", -- 0x02D8
    x"C8",x"CC",x"05",x"0F",x"90",x"EE",x"98",x"E9", -- 0x02E0
    x"08",x"8D",x"05",x"0F",x"18",x"60",x"48",x"29", -- 0x02E8
    x"DF",x"C9",x"41",x"90",x"04",x"C9",x"5B",x"90", -- 0x02F0
    x"01",x"38",x"68",x"60",x"2C",x"C7",x"10",x"30", -- 0x02F8
    x"EC",x"20",x"E1",x"83",x"20",x"C0",x"81",x"98", -- 0x0300
    x"48",x"A9",x"60",x"85",x"B0",x"A9",x"10",x"85", -- 0x0308
    x"B1",x"20",x"7E",x"83",x"A0",x"02",x"20",x"CE", -- 0x0310
    x"9F",x"20",x"35",x"83",x"20",x"35",x"83",x"20", -- 0x0318
    x"35",x"83",x"68",x"A8",x"B9",x"0E",x"0F",x"29", -- 0x0320
    x"03",x"20",x"CA",x"80",x"B9",x"0F",x"0F",x"20", -- 0x0328
    x"C2",x"80",x"4C",x"9A",x"9F",x"A2",x"03",x"B9", -- 0x0330
    x"62",x"10",x"20",x"C2",x"80",x"88",x"CA",x"D0", -- 0x0338
    x"F6",x"20",x"11",x"82",x"4C",x"CE",x"9F",x"20", -- 0x0340
    x"E1",x"83",x"4C",x"4D",x"AB",x"AD",x"CA",x"10", -- 0x0348
    x"85",x"CE",x"AD",x"CB",x"10",x"4C",x"7E",x"87", -- 0x0350
    x"20",x"BF",x"86",x"F0",x"F5",x"20",x"C5",x"FF", -- 0x0358
    x"B0",x"12",x"C9",x"3A",x"F0",x"F7",x"38",x"E9", -- 0x0360
    x"30",x"90",x"09",x"C9",x"04",x"B0",x"05",x"20", -- 0x0368
    x"7E",x"87",x"18",x"60",x"20",x"22",x"80",x"CD", -- 0x0370
    x"64",x"72",x"69",x"76",x"65",x"00",x"20",x"E1", -- 0x0378
    x"83",x"98",x"48",x"AA",x"A0",x"02",x"A9",x"00", -- 0x0380
    x"91",x"B0",x"C8",x"C0",x"12",x"D0",x"F9",x"A0", -- 0x0388
    x"02",x"20",x"CF",x"83",x"C8",x"C8",x"C0",x"0E", -- 0x0390
    x"D0",x"F7",x"68",x"AA",x"BD",x"0F",x"0E",x"10", -- 0x0398
    x"06",x"A9",x"0A",x"A0",x"0E",x"91",x"B0",x"BD", -- 0x03A0
    x"0E",x"0F",x"A0",x"04",x"20",x"BB",x"83",x"A0", -- 0x03A8
    x"0C",x"4A",x"4A",x"48",x"29",x"03",x"91",x"B0", -- 0x03B0
    x"68",x"A0",x"08",x"4A",x"4A",x"48",x"29",x"03", -- 0x03B8
    x"91",x"B0",x"C9",x"03",x"D0",x"07",x"A9",x"FF", -- 0x03C0
    x"91",x"B0",x"C8",x"91",x"B0",x"68",x"60",x"20", -- 0x03C8
    x"D2",x"83",x"BD",x"08",x"0F",x"91",x"B0",x"E8", -- 0x03D0
    x"C8",x"60",x"E6",x"AE",x"D0",x"02",x"E6",x"AF", -- 0x03D8
    x"60",x"48",x"8A",x"48",x"98",x"48",x"A9",x"84", -- 0x03E0
    x"48",x"A9",x"03",x"48",x"A0",x"05",x"BA",x"BD", -- 0x03E8
    x"07",x"01",x"48",x"88",x"D0",x"F8",x"A0",x"0A", -- 0x03F0
    x"BD",x"09",x"01",x"9D",x"0B",x"01",x"CA",x"88", -- 0x03F8
    x"D0",x"F6",x"68",x"68",x"68",x"A8",x"68",x"AA", -- 0x0400
    x"68",x"60",x"BA",x"9D",x"03",x"01",x"4C",x"04", -- 0x0408
    x"84",x"48",x"8A",x"48",x"98",x"48",x"A9",x"84", -- 0x0410
    x"48",x"A9",x"09",x"48",x"D0",x"CE",x"20",x"B8", -- 0x0418
    x"86",x"20",x"47",x"AB",x"A0",x"FF",x"84",x"A8", -- 0x0420
    x"C8",x"84",x"AA",x"B9",x"00",x"0E",x"C0",x"08", -- 0x0428
    x"90",x"03",x"B9",x"F8",x"0E",x"20",x"9C",x"80", -- 0x0430
    x"C8",x"C0",x"0C",x"D0",x"EE",x"20",x"65",x"80", -- 0x0438
    x"20",x"28",x"AD",x"04",x"0F",x"20",x"C2",x"80", -- 0x0440
    x"20",x"65",x"80",x"29",x"0D",x"44",x"72",x"69", -- 0x0448
    x"76",x"65",x"20",x"A5",x"CF",x"20",x"CA",x"80", -- 0x0450
    x"A0",x"0D",x"20",x"F4",x"81",x"20",x"65",x"80", -- 0x0458
    x"4F",x"70",x"74",x"69",x"6F",x"6E",x"20",x"AD", -- 0x0460
    x"06",x"0F",x"20",x"05",x"82",x"20",x"CA",x"80", -- 0x0468
    x"20",x"65",x"80",x"20",x"28",x"A0",x"03",x"0A", -- 0x0470
    x"0A",x"AA",x"BD",x"6F",x"85",x"20",x"9C",x"80", -- 0x0478
    x"E8",x"88",x"10",x"F6",x"20",x"65",x"80",x"29", -- 0x0480
    x"0D",x"44",x"69",x"72",x"65",x"63",x"74",x"6F", -- 0x0488
    x"72",x"79",x"20",x"3A",x"AD",x"CB",x"10",x"20", -- 0x0490
    x"CA",x"80",x"20",x"9A",x"80",x"AD",x"CA",x"10", -- 0x0498
    x"20",x"9C",x"80",x"A0",x"06",x"20",x"F4",x"81", -- 0x04A0
    x"20",x"65",x"80",x"4C",x"69",x"62",x"72",x"61", -- 0x04A8
    x"72",x"79",x"20",x"3A",x"AD",x"CD",x"10",x"20", -- 0x04B0
    x"CA",x"80",x"20",x"9A",x"80",x"AD",x"CC",x"10", -- 0x04B8
    x"20",x"9C",x"80",x"20",x"9A",x"9F",x"A0",x"00", -- 0x04C0
    x"CC",x"05",x"0F",x"B0",x"17",x"B9",x"0F",x"0E", -- 0x04C8
    x"4D",x"CA",x"10",x"29",x"7F",x"D0",x"08",x"B9", -- 0x04D0
    x"0F",x"0E",x"29",x"80",x"99",x"0F",x"0E",x"20", -- 0x04D8
    x"10",x"82",x"90",x"E4",x"A0",x"00",x"20",x"F6", -- 0x04E0
    x"84",x"90",x"16",x"A9",x"FF",x"8D",x"82",x"10", -- 0x04E8
    x"4C",x"9A",x"9F",x"20",x"10",x"82",x"CC",x"05", -- 0x04F0
    x"0F",x"B0",x"05",x"B9",x"08",x"0E",x"30",x"F3", -- 0x04F8
    x"60",x"84",x"AB",x"A2",x"00",x"B9",x"08",x"0E", -- 0x0500
    x"29",x"7F",x"9D",x"60",x"10",x"C8",x"E8",x"E0", -- 0x0508
    x"08",x"D0",x"F2",x"20",x"F6",x"84",x"B0",x"1F", -- 0x0510
    x"38",x"A2",x"06",x"B9",x"0E",x"0E",x"FD",x"60", -- 0x0518
    x"10",x"88",x"CA",x"10",x"F6",x"20",x"11",x"82", -- 0x0520
    x"B9",x"0F",x"0E",x"29",x"7F",x"ED",x"67",x"10", -- 0x0528
    x"90",x"CF",x"20",x"10",x"82",x"B0",x"DC",x"A4", -- 0x0530
    x"AB",x"B9",x"08",x"0E",x"09",x"80",x"99",x"08", -- 0x0538
    x"0E",x"AD",x"67",x"10",x"C5",x"AA",x"F0",x"10", -- 0x0540
    x"A6",x"AA",x"85",x"AA",x"D0",x"0A",x"20",x"9A", -- 0x0548
    x"9F",x"20",x"9A",x"9F",x"A0",x"FF",x"D0",x"09", -- 0x0550
    x"A4",x"A8",x"D0",x"F5",x"A0",x"05",x"20",x"F4", -- 0x0558
    x"81",x"C8",x"84",x"A8",x"A4",x"AB",x"20",x"CB", -- 0x0560
    x"9F",x"20",x"C0",x"81",x"4C",x"E4",x"84",x"6F", -- 0x0568
    x"66",x"66",x"00",x"4C",x"4F",x"41",x"44",x"52", -- 0x0570
    x"55",x"4E",x"00",x"45",x"58",x"45",x"43",x"B9", -- 0x0578
    x"0E",x"0F",x"20",x"FD",x"81",x"85",x"C4",x"18", -- 0x0580
    x"A9",x"FF",x"79",x"0C",x"0F",x"B9",x"0F",x"0F", -- 0x0588
    x"79",x"0D",x"0F",x"85",x"C5",x"B9",x"0E",x"0F", -- 0x0590
    x"29",x"03",x"65",x"C4",x"85",x"C4",x"38",x"B9", -- 0x0598
    x"07",x"0F",x"E5",x"C5",x"48",x"B9",x"06",x"0F", -- 0x05A0
    x"29",x"03",x"E5",x"C4",x"AA",x"A9",x"00",x"C5", -- 0x05A8
    x"C2",x"68",x"E5",x"C3",x"8A",x"E5",x"C6",x"60", -- 0x05B0
    x"41",x"43",x"43",x"45",x"53",x"53",x"88",x"D1", -- 0x05B8
    x"32",x"42",x"41",x"43",x"4B",x"55",x"50",x"9C", -- 0x05C0
    x"BA",x"54",x"43",x"4F",x"4D",x"50",x"41",x"43", -- 0x05C8
    x"54",x"9A",x"BF",x"0A",x"43",x"4F",x"50",x"59", -- 0x05D0
    x"9D",x"26",x"64",x"44",x"45",x"4C",x"45",x"54", -- 0x05D8
    x"45",x"86",x"FD",x"01",x"44",x"45",x"53",x"54", -- 0x05E0
    x"52",x"4F",x"59",x"87",x"0F",x"02",x"44",x"49", -- 0x05E8
    x"52",x"88",x"4D",x"09",x"44",x"52",x"49",x"56", -- 0x05F0
    x"45",x"87",x"74",x"0A",x"45",x"4E",x"41",x"42", -- 0x05F8
    x"4C",x"45",x"8A",x"38",x"00",x"49",x"4E",x"46", -- 0x0600
    x"4F",x"82",x"83",x"02",x"4C",x"49",x"42",x"88", -- 0x0608
    x"51",x"09",x"52",x"45",x"4E",x"41",x"4D",x"45", -- 0x0610
    x"8A",x"6C",x"87",x"54",x"49",x"54",x"4C",x"45", -- 0x0618
    x"88",x"A2",x"0B",x"57",x"49",x"50",x"45",x"86", -- 0x0620
    x"C2",x"02",x"B0",x"26",x"00",x"42",x"55",x"49", -- 0x0628
    x"4C",x"44",x"9F",x"47",x"01",x"43",x"41",x"52", -- 0x0630
    x"44",x"93",x"37",x"00",x"44",x"55",x"4D",x"50", -- 0x0638
    x"9E",x"CF",x"01",x"4C",x"49",x"53",x"54",x"9E", -- 0x0640
    x"8D",x"01",x"54",x"59",x"50",x"45",x"9E",x"86", -- 0x0648
    x"01",x"44",x"4D",x"4D",x"43",x"93",x"37",x"00", -- 0x0650
    x"85",x"B6",x"00",x"44",x"46",x"53",x"99",x"C5", -- 0x0658
    x"00",x"55",x"54",x"49",x"4C",x"53",x"99",x"ED", -- 0x0660
    x"00",x"99",x"F4",x"00",x"20",x"B8",x"86",x"A2", -- 0x0668
    x"FD",x"8A",x"BA",x"86",x"B6",x"AA",x"98",x"48", -- 0x0670
    x"E8",x"E8",x"68",x"48",x"A8",x"20",x"BF",x"86", -- 0x0678
    x"E8",x"BD",x"B8",x"85",x"30",x"28",x"CA",x"88", -- 0x0680
    x"86",x"B8",x"E8",x"C8",x"BD",x"B8",x"85",x"30", -- 0x0688
    x"16",x"51",x"F2",x"29",x"5F",x"F0",x"F3",x"CA", -- 0x0690
    x"E8",x"BD",x"B8",x"85",x"10",x"FA",x"B1",x"F2", -- 0x0698
    x"C9",x"2E",x"D0",x"D4",x"C8",x"B0",x"07",x"B1", -- 0x06A0
    x"F2",x"20",x"EE",x"82",x"90",x"CA",x"68",x"BD", -- 0x06A8
    x"B8",x"85",x"48",x"BD",x"B9",x"85",x"48",x"60", -- 0x06B0
    x"86",x"F2",x"84",x"F3",x"A0",x"00",x"60",x"18", -- 0x06B8
    x"4C",x"C2",x"FF",x"20",x"5E",x"82",x"20",x"01", -- 0x06C0
    x"9A",x"20",x"68",x"82",x"B9",x"0F",x"0E",x"30", -- 0x06C8
    x"12",x"20",x"C0",x"81",x"20",x"65",x"80",x"20", -- 0x06D0
    x"3A",x"20",x"EA",x"20",x"9E",x"9C",x"F0",x"09", -- 0x06D8
    x"20",x"9A",x"9F",x"20",x"9D",x"82",x"B0",x"E4", -- 0x06E0
    x"60",x"20",x"A1",x"81",x"20",x"D1",x"82",x"20", -- 0x06E8
    x"B4",x"8A",x"AC",x"CE",x"10",x"20",x"19",x"82", -- 0x06F0
    x"8C",x"CE",x"10",x"4C",x"E0",x"86",x"20",x"62", -- 0x06F8
    x"82",x"20",x"01",x"9A",x"20",x"68",x"82",x"20", -- 0x0700
    x"FC",x"82",x"20",x"D1",x"82",x"4C",x"B4",x"8A", -- 0x0708
    x"20",x"BD",x"9B",x"20",x"5E",x"82",x"20",x"01", -- 0x0710
    x"9A",x"20",x"68",x"82",x"B9",x"0F",x"0E",x"30", -- 0x0718
    x"06",x"20",x"C0",x"81",x"20",x"9A",x"9F",x"20", -- 0x0720
    x"9D",x"82",x"B0",x"F0",x"20",x"65",x"80",x"0D", -- 0x0728
    x"44",x"65",x"6C",x"65",x"74",x"65",x"20",x"28", -- 0x0730
    x"59",x"2F",x"4E",x"29",x"20",x"3F",x"20",x"EA", -- 0x0738
    x"20",x"9E",x"9C",x"F0",x"03",x"4C",x"9A",x"9F", -- 0x0740
    x"20",x"A1",x"81",x"20",x"96",x"82",x"B9",x"0F", -- 0x0748
    x"0E",x"30",x"0C",x"20",x"D1",x"82",x"AC",x"CE", -- 0x0750
    x"10",x"20",x"19",x"82",x"8C",x"CE",x"10",x"20", -- 0x0758
    x"9D",x"82",x"B0",x"EA",x"20",x"B4",x"8A",x"20", -- 0x0760
    x"65",x"80",x"0D",x"44",x"65",x"6C",x"65",x"74", -- 0x0768
    x"65",x"64",x"0D",x"EA",x"60",x"20",x"01",x"9A", -- 0x0770
    x"20",x"5D",x"83",x"8D",x"CB",x"10",x"EA",x"EA", -- 0x0778
    x"EA",x"29",x"03",x"85",x"CF",x"60",x"20",x"61", -- 0x0780
    x"89",x"20",x"6E",x"98",x"20",x"7E",x"83",x"4C", -- 0x0788
    x"A5",x"AB",x"EA",x"EA",x"20",x"6E",x"82",x"20", -- 0x0790
    x"6E",x"98",x"20",x"7E",x"83",x"84",x"BC",x"A2", -- 0x0798
    x"00",x"A5",x"C0",x"D0",x"06",x"C8",x"C8",x"A2", -- 0x07A0
    x"02",x"D0",x"08",x"B9",x"0E",x"0F",x"85",x"C4", -- 0x07A8
    x"20",x"3F",x"8A",x"B9",x"08",x"0F",x"95",x"BE", -- 0x07B0
    x"C8",x"E8",x"E0",x"08",x"D0",x"F5",x"20",x"56", -- 0x07B8
    x"8A",x"A4",x"BC",x"20",x"FC",x"82",x"4C",x"96", -- 0x07C0
    x"AB",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07C8
    x"00",x"00",x"00",x"00",x"20",x"B8",x"86",x"20", -- 0x07D0
    x"41",x"88",x"8C",x"DB",x"10",x"20",x"06",x"81", -- 0x07D8
    x"8C",x"DA",x"10",x"20",x"96",x"82",x"B0",x"22", -- 0x07E0
    x"AC",x"DB",x"10",x"AD",x"CC",x"10",x"85",x"CE", -- 0x07E8
    x"AD",x"CD",x"10",x"20",x"7E",x"87",x"20",x"09", -- 0x07F0
    x"81",x"20",x"96",x"82",x"B0",x"0C",x"20",x"22", -- 0x07F8
    x"80",x"FE",x"63",x"6F",x"6D",x"6D",x"61",x"6E", -- 0x0800
    x"64",x"00",x"20",x"9D",x"87",x"18",x"AD",x"DA", -- 0x0808
    x"10",x"A8",x"65",x"F2",x"8D",x"DA",x"10",x"A5", -- 0x0810
    x"F3",x"69",x"00",x"8D",x"DB",x"10",x"AD",x"76", -- 0x0818
    x"10",x"2D",x"77",x"10",x"0D",x"D7",x"10",x"C9", -- 0x0820
    x"FF",x"F0",x"13",x"A5",x"C0",x"8D",x"74",x"10", -- 0x0828
    x"A5",x"C1",x"8D",x"75",x"10",x"A2",x"74",x"A0", -- 0x0830
    x"10",x"A9",x"04",x"4C",x"06",x"04",x"6C",x"C0", -- 0x0838
    x"00",x"A9",x"FF",x"85",x"C0",x"A5",x"F2",x"85", -- 0x0840
    x"BC",x"A5",x"F3",x"85",x"BD",x"60",x"A2",x"00", -- 0x0848
    x"F0",x"02",x"A2",x"02",x"20",x"60",x"88",x"9D", -- 0x0850
    x"CB",x"10",x"A5",x"CE",x"9D",x"CA",x"10",x"60", -- 0x0858
    x"A9",x"24",x"85",x"CE",x"20",x"BF",x"86",x"D0", -- 0x0860
    x"07",x"A9",x"00",x"20",x"7E",x"87",x"F0",x"30", -- 0x0868
    x"AD",x"CB",x"10",x"20",x"7E",x"87",x"20",x"C5", -- 0x0870
    x"FF",x"B0",x"10",x"C9",x"3A",x"D0",x"1A",x"20", -- 0x0878
    x"5D",x"83",x"20",x"C5",x"FF",x"B0",x"19",x"C9", -- 0x0880
    x"2E",x"F0",x"EB",x"20",x"22",x"80",x"CE",x"64", -- 0x0888
    x"69",x"72",x"65",x"63",x"74",x"6F",x"72",x"79", -- 0x0890
    x"00",x"85",x"CE",x"20",x"C5",x"FF",x"90",x"EB", -- 0x0898
    x"A5",x"CF",x"60",x"20",x"01",x"9A",x"20",x"4D", -- 0x08A0
    x"83",x"20",x"47",x"83",x"4C",x"A7",x"AE",x"00", -- 0x08A8
    x"20",x"C6",x"88",x"CA",x"10",x"FA",x"E8",x"20", -- 0x08B0
    x"C5",x"FF",x"B0",x"07",x"20",x"C6",x"88",x"E0", -- 0x08B8
    x"0B",x"90",x"F3",x"4C",x"B4",x"8A",x"E0",x"08", -- 0x08C0
    x"90",x"04",x"9D",x"F8",x"0E",x"60",x"9D",x"00", -- 0x08C8
    x"0E",x"60",x"20",x"5E",x"82",x"20",x"01",x"9A", -- 0x08D0
    x"20",x"FE",x"80",x"A2",x"00",x"20",x"BF",x"86", -- 0x08D8
    x"D0",x"23",x"86",x"AA",x"20",x"96",x"82",x"B0", -- 0x08E0
    x"03",x"4C",x"76",x"82",x"20",x"4F",x"98",x"B9", -- 0x08E8
    x"0F",x"0E",x"29",x"7F",x"05",x"AA",x"99",x"0F", -- 0x08F0
    x"0E",x"20",x"FC",x"82",x"20",x"9D",x"82",x"B0", -- 0x08F8
    x"EB",x"90",x"C0",x"A2",x"80",x"20",x"C5",x"FF", -- 0x0900
    x"B0",x"D8",x"C9",x"4C",x"F0",x"F5",x"20",x"22", -- 0x0908
    x"80",x"CF",x"61",x"74",x"74",x"72",x"69",x"62", -- 0x0910
    x"75",x"74",x"65",x"00",x"20",x"E1",x"83",x"8A", -- 0x0918
    x"C9",x"04",x"F0",x"1A",x"C9",x"02",x"90",x"0B", -- 0x0920
    x"20",x"22",x"80",x"CB",x"6F",x"70",x"74",x"69", -- 0x0928
    x"6F",x"6E",x"00",x"A2",x"FF",x"98",x"F0",x"02", -- 0x0930
    x"A2",x"00",x"8E",x"C7",x"10",x"60",x"98",x"48", -- 0x0938
    x"20",x"4D",x"83",x"20",x"4D",x"AB",x"68",x"20", -- 0x0940
    x"0B",x"82",x"4D",x"06",x"0F",x"29",x"30",x"4D", -- 0x0948
    x"06",x"0F",x"8D",x"06",x"0F",x"4C",x"B4",x"8A", -- 0x0950
    x"20",x"18",x"80",x"C6",x"66",x"75",x"6C",x"6C", -- 0x0958
    x"00",x"20",x"06",x"81",x"20",x"96",x"82",x"90", -- 0x0960
    x"03",x"20",x"D1",x"82",x"A5",x"C2",x"48",x"A5", -- 0x0968
    x"C3",x"48",x"38",x"A5",x"C4",x"E5",x"C2",x"85", -- 0x0970
    x"C2",x"A5",x"C5",x"E5",x"C3",x"85",x"C3",x"AD", -- 0x0978
    x"7A",x"10",x"ED",x"78",x"10",x"85",x"C6",x"20", -- 0x0980
    x"9D",x"89",x"AD",x"79",x"10",x"8D",x"75",x"10", -- 0x0988
    x"AD",x"78",x"10",x"8D",x"74",x"10",x"68",x"85", -- 0x0990
    x"BF",x"68",x"85",x"BE",x"60",x"A9",x"00",x"85", -- 0x0998
    x"C4",x"A9",x"02",x"85",x"C5",x"AC",x"05",x"0F", -- 0x09A0
    x"F0",x"2D",x"C0",x"F8",x"B0",x"56",x"20",x"9E", -- 0x09A8
    x"85",x"4C",x"BC",x"89",x"F0",x"A2",x"20",x"19", -- 0x09B0
    x"82",x"20",x"7F",x"85",x"98",x"90",x"F5",x"84", -- 0x09B8
    x"B0",x"AC",x"05",x"0F",x"C4",x"B0",x"F0",x"0F", -- 0x09C0
    x"B9",x"07",x"0E",x"99",x"0F",x"0E",x"B9",x"07", -- 0x09C8
    x"0F",x"99",x"0F",x"0F",x"88",x"B0",x"ED",x"A2", -- 0x09D0
    x"00",x"20",x"17",x"8A",x"B5",x"C7",x"99",x"08", -- 0x09D8
    x"0E",x"C8",x"E8",x"E0",x"08",x"D0",x"F5",x"B5", -- 0x09E0
    x"BD",x"88",x"99",x"08",x"0F",x"CA",x"D0",x"F7", -- 0x09E8
    x"20",x"FC",x"82",x"98",x"48",x"AC",x"05",x"0F", -- 0x09F0
    x"20",x"10",x"82",x"8C",x"05",x"0F",x"20",x"B4", -- 0x09F8
    x"8A",x"68",x"A8",x"60",x"20",x"33",x"80",x"BE", -- 0x0A00
    x"43",x"61",x"74",x"61",x"6C",x"6F",x"67",x"75", -- 0x0A08
    x"65",x"20",x"66",x"75",x"6C",x"6C",x"00",x"AD", -- 0x0A10
    x"76",x"10",x"29",x"03",x"0A",x"0A",x"45",x"C6", -- 0x0A18
    x"29",x"FC",x"45",x"C6",x"0A",x"0A",x"4D",x"74", -- 0x0A20
    x"10",x"29",x"FC",x"4D",x"74",x"10",x"0A",x"0A", -- 0x0A28
    x"45",x"C4",x"29",x"FC",x"45",x"C4",x"85",x"C4", -- 0x0A30
    x"60",x"A9",x"01",x"8D",x"C8",x"10",x"60",x"A9", -- 0x0A38
    x"00",x"8D",x"75",x"10",x"A5",x"C4",x"20",x"FF", -- 0x0A40
    x"81",x"C9",x"03",x"D0",x"05",x"A9",x"FF",x"8D", -- 0x0A48
    x"75",x"10",x"8D",x"74",x"10",x"60",x"A9",x"00", -- 0x0A50
    x"8D",x"77",x"10",x"A5",x"C4",x"20",x"FB",x"81", -- 0x0A58
    x"C9",x"03",x"D0",x"05",x"A9",x"FF",x"8D",x"77", -- 0x0A60
    x"10",x"8D",x"76",x"10",x"60",x"20",x"62",x"82", -- 0x0A68
    x"20",x"BF",x"86",x"D0",x"03",x"4C",x"06",x"9A", -- 0x0A70
    x"20",x"FE",x"80",x"98",x"48",x"20",x"96",x"82", -- 0x0A78
    x"B0",x"03",x"4C",x"76",x"82",x"20",x"4C",x"98", -- 0x0A80
    x"84",x"B3",x"68",x"A8",x"20",x"BF",x"86",x"F0", -- 0x0A88
    x"E4",x"20",x"FE",x"80",x"20",x"96",x"82",x"90", -- 0x0A90
    x"0B",x"20",x"2B",x"80",x"C4",x"65",x"78",x"69", -- 0x0A98
    x"73",x"74",x"73",x"00",x"A4",x"B3",x"20",x"10", -- 0x0AA0
    x"82",x"A2",x"07",x"B5",x"C7",x"99",x"07",x"0E", -- 0x0AA8
    x"88",x"CA",x"10",x"F7",x"18",x"F8",x"AD",x"04", -- 0x0AB0
    x"0F",x"69",x"01",x"D8",x"8D",x"04",x"0F",x"4C", -- 0x0AB8
    x"61",x"AB",x"A9",x"FF",x"20",x"9E",x"06",x"AD", -- 0x0AC0
    x"E3",x"FE",x"A9",x"00",x"20",x"95",x"06",x"A8", -- 0x0AC8
    x"B1",x"FD",x"20",x"95",x"06",x"C8",x"B1",x"FD", -- 0x0AD0
    x"20",x"95",x"06",x"AA",x"D0",x"F7",x"A2",x"FF", -- 0x0AD8
    x"9A",x"58",x"2C",x"E0",x"FE",x"10",x"06",x"AD", -- 0x0AE0
    x"E1",x"FE",x"20",x"EE",x"FF",x"2C",x"E2",x"FE", -- 0x0AE8
    x"10",x"F0",x"2C",x"E0",x"FE",x"30",x"F0",x"AE", -- 0x0AF0
    x"E3",x"FE",x"86",x"51",x"6C",x"00",x"05",x"00", -- 0x0AF8
    x"80",x"00",x"00",x"4C",x"84",x"04",x"4C",x"A7", -- 0x0B00
    x"06",x"C9",x"80",x"90",x"2B",x"C9",x"C0",x"B0", -- 0x0B08
    x"1A",x"09",x"40",x"C5",x"15",x"D0",x"20",x"08", -- 0x0B10
    x"78",x"A9",x"05",x"20",x"9E",x"06",x"A5",x"15", -- 0x0B18
    x"20",x"9E",x"06",x"28",x"A9",x"80",x"85",x"15", -- 0x0B20
    x"85",x"14",x"60",x"06",x"14",x"B0",x"06",x"C5", -- 0x0B28
    x"15",x"F0",x"04",x"18",x"60",x"85",x"15",x"60", -- 0x0B30
    x"08",x"78",x"84",x"13",x"86",x"12",x"20",x"9E", -- 0x0B38
    x"06",x"AA",x"A0",x"03",x"A5",x"15",x"20",x"9E", -- 0x0B40
    x"06",x"B1",x"12",x"20",x"9E",x"06",x"88",x"10", -- 0x0B48
    x"F8",x"A0",x"18",x"8C",x"E0",x"FE",x"BD",x"18", -- 0x0B50
    x"05",x"8D",x"E0",x"FE",x"4A",x"4A",x"90",x"06", -- 0x0B58
    x"2C",x"E5",x"FE",x"2C",x"E5",x"FE",x"20",x"9E", -- 0x0B60
    x"06",x"2C",x"E6",x"FE",x"50",x"FB",x"B0",x"0D", -- 0x0B68
    x"E0",x"04",x"D0",x"11",x"20",x"14",x"04",x"20", -- 0x0B70
    x"95",x"06",x"4C",x"32",x"00",x"4A",x"90",x"05", -- 0x0B78
    x"A0",x"88",x"8C",x"E0",x"FE",x"28",x"60",x"58", -- 0x0B80
    x"B0",x"11",x"D0",x"03",x"4C",x"9C",x"05",x"A2", -- 0x0B88
    x"00",x"A0",x"FF",x"A9",x"FD",x"20",x"F4",x"FF", -- 0x0B90
    x"8A",x"F0",x"D9",x"A9",x"FF",x"20",x"06",x"04", -- 0x0B98
    x"90",x"F9",x"20",x"D2",x"04",x"A9",x"07",x"20", -- 0x0BA0
    x"CB",x"04",x"A0",x"00",x"84",x"00",x"B1",x"00", -- 0x0BA8
    x"8D",x"E5",x"FE",x"EA",x"EA",x"EA",x"C8",x"D0", -- 0x0BB0
    x"F5",x"E6",x"54",x"D0",x"06",x"E6",x"55",x"D0", -- 0x0BB8
    x"02",x"E6",x"56",x"E6",x"01",x"24",x"01",x"50", -- 0x0BC0
    x"DC",x"20",x"D2",x"04",x"A9",x"04",x"A0",x"00", -- 0x0BC8
    x"A2",x"53",x"4C",x"06",x"04",x"A9",x"80",x"85", -- 0x0BD0
    x"54",x"85",x"01",x"A9",x"20",x"2D",x"06",x"80", -- 0x0BD8
    x"A8",x"84",x"53",x"F0",x"19",x"AE",x"07",x"80", -- 0x0BE0
    x"E8",x"BD",x"00",x"80",x"D0",x"FA",x"BD",x"01", -- 0x0BE8
    x"80",x"85",x"53",x"BD",x"02",x"80",x"85",x"54", -- 0x0BF0
    x"BC",x"03",x"80",x"BD",x"04",x"80",x"85",x"56", -- 0x0BF8
    x"84",x"55",x"60",x"37",x"05",x"96",x"05",x"F2", -- 0x0C00
    x"05",x"07",x"06",x"27",x"06",x"68",x"06",x"5E", -- 0x0C08
    x"05",x"2D",x"05",x"20",x"05",x"42",x"05",x"A9", -- 0x0C10
    x"05",x"D1",x"05",x"86",x"88",x"96",x"98",x"18", -- 0x0C18
    x"18",x"82",x"18",x"20",x"C5",x"06",x"A8",x"20", -- 0x0C20
    x"C5",x"06",x"20",x"D4",x"FF",x"4C",x"9C",x"05", -- 0x0C28
    x"20",x"C5",x"06",x"A8",x"20",x"D7",x"FF",x"4C", -- 0x0C30
    x"3A",x"05",x"20",x"E0",x"FF",x"6A",x"20",x"95", -- 0x0C38
    x"06",x"2A",x"4C",x"9E",x"05",x"20",x"C5",x"06", -- 0x0C40
    x"F0",x"0B",x"48",x"20",x"82",x"05",x"68",x"20", -- 0x0C48
    x"CE",x"FF",x"4C",x"9E",x"05",x"20",x"C5",x"06", -- 0x0C50
    x"A8",x"A9",x"00",x"20",x"CE",x"FF",x"4C",x"9C", -- 0x0C58
    x"05",x"20",x"C5",x"06",x"A8",x"A2",x"04",x"20", -- 0x0C60
    x"C5",x"06",x"95",x"FF",x"CA",x"D0",x"F8",x"20", -- 0x0C68
    x"C5",x"06",x"20",x"DA",x"FF",x"20",x"95",x"06", -- 0x0C70
    x"A2",x"03",x"B5",x"00",x"20",x"95",x"06",x"CA", -- 0x0C78
    x"10",x"F8",x"4C",x"36",x"00",x"A2",x"00",x"A0", -- 0x0C80
    x"00",x"20",x"C5",x"06",x"99",x"00",x"07",x"C8", -- 0x0C88
    x"F0",x"04",x"C9",x"0D",x"D0",x"F3",x"A0",x"07", -- 0x0C90
    x"60",x"20",x"82",x"05",x"20",x"F7",x"FF",x"A9", -- 0x0C98
    x"7F",x"2C",x"E2",x"FE",x"50",x"FB",x"8D",x"E3", -- 0x0CA0
    x"FE",x"4C",x"36",x"00",x"A2",x"10",x"20",x"C5", -- 0x0CA8
    x"06",x"95",x"01",x"CA",x"D0",x"F8",x"20",x"82", -- 0x0CB0
    x"05",x"86",x"00",x"84",x"01",x"A0",x"00",x"20", -- 0x0CB8
    x"C5",x"06",x"20",x"DD",x"FF",x"20",x"95",x"06", -- 0x0CC0
    x"A2",x"10",x"B5",x"01",x"20",x"95",x"06",x"CA", -- 0x0CC8
    x"D0",x"F8",x"F0",x"D5",x"A2",x"0D",x"20",x"C5", -- 0x0CD0
    x"06",x"95",x"FF",x"CA",x"D0",x"F8",x"20",x"C5", -- 0x0CD8
    x"06",x"A0",x"00",x"20",x"D1",x"FF",x"48",x"A2", -- 0x0CE0
    x"0C",x"B5",x"00",x"20",x"95",x"06",x"CA",x"10", -- 0x0CE8
    x"F8",x"68",x"4C",x"3A",x"05",x"20",x"C5",x"06", -- 0x0CF0
    x"AA",x"20",x"C5",x"06",x"20",x"F4",x"FF",x"2C", -- 0x0CF8
    x"E2",x"FE",x"50",x"FB",x"8E",x"E3",x"FE",x"4C", -- 0x0D00
    x"36",x"00",x"20",x"C5",x"06",x"AA",x"20",x"C5", -- 0x0D08
    x"06",x"A8",x"20",x"C5",x"06",x"20",x"F4",x"FF", -- 0x0D10
    x"49",x"9D",x"F0",x"EB",x"6A",x"20",x"95",x"06", -- 0x0D18
    x"2C",x"E2",x"FE",x"50",x"FB",x"8C",x"E3",x"FE", -- 0x0D20
    x"70",x"D5",x"20",x"C5",x"06",x"A8",x"2C",x"E2", -- 0x0D28
    x"FE",x"10",x"FB",x"AE",x"E3",x"FE",x"CA",x"30", -- 0x0D30
    x"0F",x"2C",x"E2",x"FE",x"10",x"FB",x"AD",x"E3", -- 0x0D38
    x"FE",x"9D",x"28",x"01",x"CA",x"10",x"F2",x"98", -- 0x0D40
    x"A2",x"28",x"A0",x"01",x"20",x"F1",x"FF",x"2C", -- 0x0D48
    x"E2",x"FE",x"10",x"FB",x"AE",x"E3",x"FE",x"CA", -- 0x0D50
    x"30",x"0E",x"BC",x"28",x"01",x"2C",x"E2",x"FE", -- 0x0D58
    x"50",x"FB",x"8C",x"E3",x"FE",x"CA",x"10",x"F2", -- 0x0D60
    x"4C",x"36",x"00",x"A2",x"04",x"20",x"C5",x"06", -- 0x0D68
    x"95",x"00",x"CA",x"10",x"F8",x"E8",x"A0",x"00", -- 0x0D70
    x"8A",x"20",x"F1",x"FF",x"90",x"05",x"A9",x"FF", -- 0x0D78
    x"4C",x"9E",x"05",x"A2",x"00",x"A9",x"7F",x"20", -- 0x0D80
    x"95",x"06",x"BD",x"00",x"07",x"20",x"95",x"06", -- 0x0D88
    x"E8",x"C9",x"0D",x"D0",x"F5",x"4C",x"36",x"00", -- 0x0D90
    x"2C",x"E2",x"FE",x"50",x"FB",x"8D",x"E3",x"FE", -- 0x0D98
    x"60",x"2C",x"E6",x"FE",x"50",x"FB",x"8D",x"E7", -- 0x0DA0
    x"FE",x"60",x"A5",x"FF",x"38",x"6A",x"30",x"0F", -- 0x0DA8
    x"48",x"A9",x"00",x"20",x"BC",x"06",x"98",x"20", -- 0x0DB0
    x"BC",x"06",x"8A",x"20",x"BC",x"06",x"68",x"2C", -- 0x0DB8
    x"E0",x"FE",x"50",x"FB",x"8D",x"E1",x"FE",x"60", -- 0x0DC0
    x"2C",x"E2",x"FE",x"10",x"FB",x"AD",x"E3",x"FE", -- 0x0DC8
    x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DD0
    x"00",x"00",x"00",x"00",x"00",x"A2",x"11",x"A0", -- 0x0DD8
    x"15",x"60",x"20",x"E1",x"83",x"A9",x"77",x"4C", -- 0x0DE0
    x"F4",x"FF",x"20",x"E2",x"8D",x"A9",x"00",x"18", -- 0x0DE8
    x"69",x"20",x"F0",x"ED",x"A8",x"20",x"05",x"8E", -- 0x0DF0
    x"D0",x"F5",x"98",x"F0",x"ED",x"20",x"7B",x"90", -- 0x0DF8
    x"90",x"03",x"4C",x"AD",x"90",x"48",x"20",x"51", -- 0x0E00
    x"90",x"B0",x"45",x"B9",x"1B",x"11",x"49",x"FF", -- 0x0E08
    x"2D",x"C0",x"10",x"8D",x"C0",x"10",x"B9",x"17", -- 0x0E10
    x"11",x"29",x"60",x"F0",x"33",x"20",x"55",x"8E", -- 0x0E18
    x"B9",x"17",x"11",x"29",x"20",x"F0",x"26",x"AE", -- 0x0E20
    x"C4",x"10",x"B9",x"14",x"11",x"9D",x"0C",x"0F", -- 0x0E28
    x"B9",x"15",x"11",x"9D",x"0D",x"0F",x"B9",x"16", -- 0x0E30
    x"11",x"20",x"0B",x"82",x"5D",x"0E",x"0F",x"29", -- 0x0E38
    x"30",x"5D",x"0E",x"0F",x"9D",x"0E",x"0F",x"20", -- 0x0E40
    x"B4",x"8A",x"AC",x"C2",x"10",x"20",x"4B",x"91", -- 0x0E48
    x"AE",x"C6",x"10",x"68",x"60",x"20",x"83",x"8E", -- 0x0E50
    x"A2",x"07",x"B9",x"0C",x"11",x"95",x"C6",x"88", -- 0x0E58
    x"88",x"CA",x"D0",x"F6",x"20",x"96",x"82",x"90", -- 0x0E60
    x"27",x"8C",x"C4",x"10",x"B9",x"0E",x"0F",x"BE", -- 0x0E68
    x"0F",x"0F",x"AC",x"C2",x"10",x"59",x"0D",x"11", -- 0x0E70
    x"29",x"03",x"D0",x"14",x"8A",x"D9",x"0F",x"11", -- 0x0E78
    x"D0",x"0E",x"60",x"B9",x"0E",x"11",x"29",x"7F", -- 0x0E80
    x"85",x"CE",x"B9",x"17",x"11",x"4C",x"7E",x"87", -- 0x0E88
    x"4C",x"AF",x"81",x"C9",x"00",x"D0",x"06",x"20", -- 0x0E90
    x"E1",x"83",x"4C",x"FA",x"8D",x"20",x"11",x"84", -- 0x0E98
    x"86",x"BC",x"84",x"BD",x"85",x"B4",x"24",x"B4", -- 0x0EA0
    x"08",x"20",x"06",x"81",x"20",x"96",x"82",x"B0", -- 0x0EA8
    x"1A",x"28",x"50",x"03",x"A9",x"00",x"60",x"08", -- 0x0EB0
    x"A9",x"00",x"A2",x"07",x"95",x"BE",x"9D",x"74", -- 0x0EB8
    x"10",x"CA",x"10",x"F8",x"A9",x"40",x"85",x"C5", -- 0x0EC0
    x"20",x"61",x"89",x"28",x"08",x"70",x"03",x"20", -- 0x0EC8
    x"3C",x"98",x"20",x"9E",x"8F",x"90",x"0E",x"B9", -- 0x0ED0
    x"0C",x"11",x"10",x"26",x"24",x"B4",x"30",x"22", -- 0x0ED8
    x"20",x"99",x"8F",x"B0",x"F2",x"AC",x"C2",x"10", -- 0x0EE0
    x"D0",x"21",x"20",x"33",x"80",x"C0",x"54",x"6F", -- 0x0EE8
    x"6F",x"20",x"6D",x"61",x"6E",x"79",x"20",x"66", -- 0x0EF0
    x"69",x"6C",x"65",x"73",x"20",x"6F",x"70",x"65", -- 0x0EF8
    x"6E",x"00",x"20",x"2B",x"80",x"C2",x"6F",x"70", -- 0x0F00
    x"65",x"6E",x"00",x"A9",x"08",x"8D",x"C5",x"10", -- 0x0F08
    x"BD",x"08",x"0E",x"99",x"00",x"11",x"C8",x"BD", -- 0x0F10
    x"08",x"0F",x"99",x"00",x"11",x"C8",x"E8",x"CE", -- 0x0F18
    x"C5",x"10",x"D0",x"EC",x"A2",x"10",x"A9",x"00", -- 0x0F20
    x"99",x"00",x"11",x"C8",x"CA",x"D0",x"F9",x"AD", -- 0x0F28
    x"C2",x"10",x"A8",x"20",x"04",x"82",x"69",x"11", -- 0x0F30
    x"99",x"13",x"11",x"AD",x"C1",x"10",x"99",x"1B", -- 0x0F38
    x"11",x"0D",x"C0",x"10",x"8D",x"C0",x"10",x"B9", -- 0x0F40
    x"09",x"11",x"69",x"FF",x"B9",x"0B",x"11",x"69", -- 0x0F48
    x"00",x"99",x"19",x"11",x"B9",x"0D",x"11",x"09", -- 0x0F50
    x"0F",x"69",x"00",x"20",x"FD",x"81",x"99",x"1A", -- 0x0F58
    x"11",x"28",x"50",x"2E",x"30",x"08",x"A9",x"80", -- 0x0F60
    x"19",x"0C",x"11",x"99",x"0C",x"11",x"B9",x"09", -- 0x0F68
    x"11",x"99",x"14",x"11",x"B9",x"0B",x"11",x"99", -- 0x0F70
    x"15",x"11",x"B9",x"0D",x"11",x"20",x"FD",x"81", -- 0x0F78
    x"99",x"16",x"11",x"A5",x"CF",x"19",x"17",x"11", -- 0x0F80
    x"99",x"17",x"11",x"98",x"20",x"04",x"82",x"09", -- 0x0F88
    x"10",x"60",x"A9",x"20",x"99",x"17",x"11",x"D0", -- 0x0F90
    x"EA",x"8A",x"48",x"4C",x"DD",x"8F",x"A9",x"00", -- 0x0F98
    x"8D",x"C2",x"10",x"A9",x"08",x"85",x"B5",x"98", -- 0x0FA0
    x"AA",x"A0",x"A0",x"84",x"B3",x"8A",x"48",x"A9", -- 0x0FA8
    x"08",x"85",x"B2",x"A5",x"B5",x"2C",x"C0",x"10", -- 0x0FB0
    x"F0",x"1D",x"B9",x"17",x"11",x"45",x"CF",x"29", -- 0x0FB8
    x"03",x"D0",x"1A",x"BD",x"08",x"0E",x"59",x"00", -- 0x0FC0
    x"11",x"29",x"7F",x"D0",x"10",x"E8",x"C8",x"C8", -- 0x0FC8
    x"C6",x"B2",x"D0",x"EF",x"38",x"B0",x"10",x"8C", -- 0x0FD0
    x"C2",x"10",x"8D",x"C1",x"10",x"38",x"A5",x"B3", -- 0x0FD8
    x"E9",x"20",x"85",x"B3",x"06",x"B5",x"18",x"68", -- 0x0FE0
    x"AA",x"A4",x"B3",x"A5",x"B5",x"B0",x"02",x"D0", -- 0x0FE8
    x"BA",x"60",x"AD",x"C0",x"10",x"48",x"20",x"ED", -- 0x0FF0
    x"8D",x"F0",x"07",x"AD",x"C0",x"10",x"48",x"20", -- 0x0FF8
    x"FA",x"8D",x"68",x"8D",x"C0",x"10",x"60",x"C0", -- 0x1000
    x"00",x"F0",x"11",x"20",x"E1",x"83",x"C9",x"FF", -- 0x1008
    x"F0",x"E9",x"C9",x"03",x"B0",x"17",x"4A",x"90", -- 0x1010
    x"15",x"4C",x"A7",x"92",x"20",x"11",x"84",x"A8", -- 0x1018
    x"C8",x"C0",x"03",x"B0",x"08",x"B9",x"81",x"99", -- 0x1020
    x"48",x"B9",x"7E",x"99",x"48",x"60",x"20",x"E1", -- 0x1028
    x"83",x"20",x"A5",x"90",x"8C",x"C2",x"10",x"0A", -- 0x1030
    x"0A",x"6D",x"C2",x"10",x"A8",x"B9",x"10",x"11", -- 0x1038
    x"95",x"00",x"B9",x"11",x"11",x"95",x"01",x"B9", -- 0x1040
    x"12",x"11",x"95",x"02",x"A9",x"00",x"95",x"03", -- 0x1048
    x"60",x"48",x"8E",x"C6",x"10",x"98",x"29",x"E0", -- 0x1050
    x"8D",x"C2",x"10",x"F0",x"13",x"20",x"04",x"82", -- 0x1058
    x"A8",x"A9",x"00",x"38",x"6A",x"88",x"D0",x"FC", -- 0x1060
    x"AC",x"C2",x"10",x"2C",x"C0",x"10",x"D0",x"03", -- 0x1068
    x"68",x"38",x"60",x"68",x"18",x"60",x"48",x"8A", -- 0x1070
    x"4C",x"7D",x"90",x"48",x"98",x"C9",x"10",x"90", -- 0x1078
    x"04",x"C9",x"18",x"90",x"02",x"A9",x"08",x"20", -- 0x1080
    x"0A",x"82",x"A8",x"68",x"60",x"48",x"98",x"48", -- 0x1088
    x"8A",x"A8",x"20",x"A5",x"90",x"98",x"20",x"F8", -- 0x1090
    x"92",x"D0",x"04",x"A2",x"FF",x"D0",x"02",x"A2", -- 0x1098
    x"00",x"68",x"A8",x"68",x"60",x"20",x"7B",x"90", -- 0x10A0
    x"20",x"51",x"90",x"90",x"F7",x"20",x"33",x"80", -- 0x10A8
    x"DE",x"43",x"68",x"61",x"6E",x"6E",x"65",x"6C", -- 0x10B0
    x"00",x"20",x"33",x"80",x"DF",x"45",x"4F",x"46", -- 0x10B8
    x"00",x"20",x"11",x"84",x"20",x"A5",x"90",x"98", -- 0x10C0
    x"20",x"F8",x"92",x"D0",x"13",x"B9",x"17",x"11", -- 0x10C8
    x"29",x"10",x"D0",x"E5",x"A9",x"10",x"20",x"3C", -- 0x10D0
    x"91",x"AE",x"C6",x"10",x"A9",x"FE",x"38",x"60", -- 0x10D8
    x"B9",x"17",x"11",x"30",x"0A",x"20",x"83",x"8E", -- 0x10E0
    x"20",x"4B",x"91",x"38",x"20",x"53",x"91",x"B9", -- 0x10E8
    x"10",x"11",x"85",x"BC",x"B9",x"13",x"11",x"85", -- 0x10F0
    x"BD",x"A0",x"00",x"B1",x"BC",x"48",x"AC",x"C2", -- 0x10F8
    x"10",x"A6",x"BC",x"E8",x"8A",x"99",x"10",x"11", -- 0x1100
    x"D0",x"14",x"18",x"B9",x"11",x"11",x"69",x"01", -- 0x1108
    x"99",x"11",x"11",x"B9",x"12",x"11",x"69",x"00", -- 0x1110
    x"99",x"12",x"11",x"20",x"41",x"91",x"18",x"68", -- 0x1118
    x"60",x"18",x"B9",x"0F",x"11",x"79",x"11",x"11", -- 0x1120
    x"85",x"C5",x"99",x"1C",x"11",x"B9",x"0D",x"11", -- 0x1128
    x"29",x"03",x"79",x"12",x"11",x"85",x"C4",x"99", -- 0x1130
    x"1D",x"11",x"A9",x"80",x"19",x"17",x"11",x"D0", -- 0x1138
    x"05",x"A9",x"7F",x"39",x"17",x"11",x"99",x"17", -- 0x1140
    x"11",x"18",x"60",x"B9",x"17",x"11",x"29",x"40", -- 0x1148
    x"F0",x"3D",x"18",x"08",x"20",x"0B",x"B9",x"AC", -- 0x1150
    x"C2",x"10",x"B9",x"13",x"11",x"85",x"BF",x"20", -- 0x1158
    x"8D",x"A0",x"A9",x"00",x"85",x"BE",x"85",x"C2", -- 0x1160
    x"A9",x"01",x"85",x"C3",x"28",x"B0",x"17",x"B9", -- 0x1168
    x"1C",x"11",x"85",x"C5",x"B9",x"1D",x"11",x"85", -- 0x1170
    x"C4",x"20",x"8F",x"87",x"AC",x"C2",x"10",x"A9", -- 0x1178
    x"BF",x"20",x"43",x"91",x"90",x"06",x"20",x"21", -- 0x1180
    x"91",x"20",x"C6",x"87",x"AC",x"C2",x"10",x"60", -- 0x1188
    x"4C",x"AD",x"90",x"4C",x"41",x"98",x"20",x"2B", -- 0x1190
    x"80",x"C1",x"72",x"65",x"61",x"64",x"20",x"6F", -- 0x1198
    x"6E",x"6C",x"79",x"00",x"20",x"E1",x"83",x"4C", -- 0x11A0
    x"B0",x"91",x"20",x"E1",x"83",x"20",x"A5",x"90", -- 0x11A8
    x"48",x"B9",x"0C",x"11",x"30",x"E0",x"B9",x"0E", -- 0x11B0
    x"11",x"30",x"D8",x"20",x"83",x"8E",x"98",x"18", -- 0x11B8
    x"69",x"04",x"20",x"F8",x"92",x"D0",x"76",x"20", -- 0x11C0
    x"58",x"8E",x"AE",x"C4",x"10",x"38",x"BD",x"07", -- 0x11C8
    x"0F",x"FD",x"0F",x"0F",x"48",x"BD",x"06",x"0F", -- 0x11D0
    x"FD",x"0E",x"0F",x"29",x"03",x"8D",x"C3",x"10", -- 0x11D8
    x"0A",x"0A",x"0A",x"0A",x"5D",x"0E",x"0F",x"29", -- 0x11E0
    x"30",x"5D",x"0E",x"0F",x"9D",x"0E",x"0F",x"AD", -- 0x11E8
    x"C3",x"10",x"D9",x"1A",x"11",x"D0",x"2B",x"68", -- 0x11F0
    x"D9",x"19",x"11",x"D0",x"26",x"84",x"B4",x"20", -- 0x11F8
    x"20",x"99",x"20",x"76",x"90",x"C4",x"B4",x"D0", -- 0x1200
    x"03",x"20",x"11",x"99",x"A4",x"B4",x"20",x"05", -- 0x1208
    x"8E",x"20",x"33",x"80",x"BF",x"43",x"61",x"6E", -- 0x1210
    x"27",x"74",x"20",x"65",x"78",x"74",x"65",x"6E", -- 0x1218
    x"64",x"00",x"68",x"9D",x"0D",x"0F",x"99",x"19", -- 0x1220
    x"11",x"AD",x"C3",x"10",x"99",x"1A",x"11",x"A9", -- 0x1228
    x"00",x"9D",x"0C",x"0F",x"20",x"B4",x"8A",x"EA", -- 0x1230
    x"EA",x"EA",x"AC",x"C2",x"10",x"B9",x"17",x"11", -- 0x1238
    x"30",x"17",x"20",x"4B",x"91",x"B9",x"14",x"11", -- 0x1240
    x"D0",x"0B",x"98",x"20",x"F8",x"92",x"D0",x"05", -- 0x1248
    x"20",x"21",x"91",x"D0",x"04",x"38",x"20",x"53", -- 0x1250
    x"91",x"B9",x"10",x"11",x"85",x"BC",x"B9",x"13", -- 0x1258
    x"11",x"85",x"BD",x"68",x"A0",x"00",x"91",x"BC", -- 0x1260
    x"AC",x"C2",x"10",x"A9",x"40",x"20",x"3C",x"91", -- 0x1268
    x"E6",x"BC",x"A5",x"BC",x"99",x"10",x"11",x"D0", -- 0x1270
    x"13",x"20",x"41",x"91",x"B9",x"11",x"11",x"69", -- 0x1278
    x"01",x"99",x"11",x"11",x"B9",x"12",x"11",x"69", -- 0x1280
    x"00",x"99",x"12",x"11",x"98",x"20",x"F8",x"92", -- 0x1288
    x"90",x"14",x"A9",x"20",x"20",x"3C",x"91",x"A2", -- 0x1290
    x"02",x"B9",x"10",x"11",x"99",x"14",x"11",x"C8", -- 0x1298
    x"CA",x"10",x"F6",x"88",x"88",x"88",x"60",x"20", -- 0x12A0
    x"E1",x"83",x"20",x"A5",x"90",x"20",x"5E",x"A1", -- 0x12A8
    x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"20",x"10", -- 0x12B0
    x"93",x"B0",x"08",x"A9",x"00",x"20",x"A4",x"91", -- 0x12B8
    x"4C",x"B6",x"92",x"B5",x"00",x"99",x"10",x"11", -- 0x12C0
    x"B5",x"01",x"99",x"11",x"11",x"B5",x"02",x"99", -- 0x12C8
    x"12",x"11",x"A9",x"6F",x"20",x"43",x"91",x"B9", -- 0x12D0
    x"0F",x"11",x"79",x"11",x"11",x"8D",x"C5",x"10", -- 0x12D8
    x"B9",x"0D",x"11",x"29",x"03",x"79",x"12",x"11", -- 0x12E0
    x"D9",x"1D",x"11",x"D0",x"B9",x"AD",x"C5",x"10", -- 0x12E8
    x"D9",x"1C",x"11",x"D0",x"B1",x"4C",x"3A",x"91", -- 0x12F0
    x"AA",x"B9",x"12",x"11",x"DD",x"16",x"11",x"D0", -- 0x12F8
    x"0E",x"B9",x"11",x"11",x"DD",x"15",x"11",x"D0", -- 0x1300
    x"06",x"B9",x"10",x"11",x"DD",x"14",x"11",x"60", -- 0x1308
    x"B9",x"14",x"11",x"D5",x"00",x"B9",x"15",x"11", -- 0x1310
    x"F5",x"01",x"B9",x"16",x"11",x"F5",x"02",x"60", -- 0x1318
    x"A5",x"B3",x"48",x"A9",x"FF",x"8D",x"DE",x"10", -- 0x1320
    x"20",x"65",x"80",x"53",x"75",x"70",x"65",x"72", -- 0x1328
    x"20",x"4D",x"4D",x"43",x"0D",x"0D",x"90",x"03", -- 0x1330
    x"4C",x"55",x"A1",x"A9",x"00",x"BA",x"9D",x"06", -- 0x1338
    x"01",x"A9",x"06",x"20",x"15",x"80",x"A2",x"0D", -- 0x1340
    x"BD",x"49",x"99",x"9D",x"12",x"02",x"CA",x"10", -- 0x1348
    x"F7",x"20",x"28",x"99",x"84",x"B1",x"86",x"B0", -- 0x1350
    x"A2",x"07",x"A0",x"1B",x"B9",x"3C",x"99",x"91", -- 0x1358
    x"B0",x"C8",x"B9",x"3C",x"99",x"91",x"B0",x"C8", -- 0x1360
    x"A5",x"F4",x"91",x"B0",x"C8",x"CA",x"D0",x"EC", -- 0x1368
    x"86",x"CF",x"8C",x"82",x"10",x"A2",x"0F",x"20", -- 0x1370
    x"2C",x"99",x"20",x"9E",x"98",x"A0",x"D4",x"B1", -- 0x1378
    x"B0",x"10",x"2F",x"A0",x"D5",x"B1",x"B0",x"30", -- 0x1380
    x"27",x"20",x"8F",x"98",x"A0",x"00",x"B1",x"B0", -- 0x1388
    x"C0",x"C0",x"90",x"05",x"99",x"00",x"10",x"B0", -- 0x1390
    x"03",x"99",x"00",x"11",x"88",x"D0",x"EF",x"A9", -- 0x1398
    x"A0",x"A8",x"48",x"A9",x"3F",x"20",x"43",x"91", -- 0x13A0
    x"68",x"99",x"1D",x"11",x"E9",x"1F",x"D0",x"F1", -- 0x13A8
    x"68",x"60",x"A9",x"FF",x"91",x"B0",x"8D",x"D4", -- 0x13B0
    x"10",x"20",x"8F",x"98",x"20",x"24",x"99",x"8A", -- 0x13B8
    x"49",x"FF",x"8D",x"D7",x"10",x"A9",x"24",x"8D", -- 0x13C0
    x"CA",x"10",x"8D",x"CC",x"10",x"A0",x"00",x"8C", -- 0x13C8
    x"CB",x"10",x"8C",x"CD",x"10",x"A0",x"00",x"8C", -- 0x13D0
    x"C0",x"10",x"8C",x"C9",x"10",x"88",x"8C",x"C8", -- 0x13D8
    x"10",x"8C",x"C7",x"10",x"8C",x"DE",x"10",x"20", -- 0x13E0
    x"0A",x"AD",x"4C",x"04",x"94",x"00",x"00",x"00", -- 0x13E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x13F8
    x"00",x"00",x"00",x"00",x"68",x"D0",x"34",x"20", -- 0x1400
    x"4D",x"AB",x"A0",x"00",x"A2",x"00",x"AD",x"06", -- 0x1408
    x"0F",x"20",x"05",x"82",x"F0",x"25",x"48",x"A2", -- 0x1410
    x"43",x"A0",x"99",x"20",x"B8",x"86",x"20",x"FE", -- 0x1418
    x"80",x"20",x"96",x"82",x"68",x"B0",x"15",x"20", -- 0x1420
    x"65",x"80",x"46",x"69",x"6C",x"65",x"20",x"6E", -- 0x1428
    x"6F",x"74",x"20",x"66",x"6F",x"75",x"6E",x"64", -- 0x1430
    x"0D",x"0D",x"EA",x"60",x"C9",x"02",x"90",x"0E", -- 0x1438
    x"F0",x"06",x"A2",x"41",x"A0",x"99",x"D0",x"0A", -- 0x1440
    x"A2",x"43",x"A0",x"99",x"D0",x"04",x"A2",x"39", -- 0x1448
    x"A0",x"99",x"4C",x"F7",x"FF",x"C9",x"01",x"D0", -- 0x1450
    x"07",x"C0",x"17",x"B0",x"02",x"A0",x"17",x"60", -- 0x1458
    x"C9",x"02",x"D0",x"1A",x"48",x"98",x"18",x"85", -- 0x1460
    x"B1",x"9D",x"F0",x"0D",x"69",x"02",x"48",x"A9", -- 0x1468
    x"00",x"85",x"B0",x"A0",x"D4",x"91",x"B0",x"C8", -- 0x1470
    x"91",x"B0",x"68",x"A8",x"68",x"60",x"C9",x"03", -- 0x1478
    x"D0",x"19",x"84",x"B3",x"20",x"E1",x"83",x"4C", -- 0x1480
    x"F7",x"A7",x"F4",x"FF",x"8A",x"30",x"09",x"C9", -- 0x1488
    x"32",x"D0",x"EA",x"A9",x"78",x"20",x"F4",x"FF", -- 0x1490
    x"4C",x"20",x"93",x"C9",x"04",x"D0",x"08",x"20", -- 0x1498
    x"E1",x"83",x"A2",x"72",x"4C",x"71",x"86",x"C9", -- 0x14A0
    x"09",x"D0",x"12",x"20",x"E1",x"83",x"4C",x"94", -- 0x14A8
    x"AF",x"A0",x"C9",x"0D",x"D0",x"EE",x"98",x"E8", -- 0x14B0
    x"A0",x"02",x"4C",x"CB",x"99",x"C9",x"0A",x"D0", -- 0x14B8
    x"29",x"20",x"E1",x"83",x"20",x"9E",x"98",x"A0", -- 0x14C0
    x"D5",x"B1",x"B0",x"10",x"1C",x"A0",x"00",x"C0", -- 0x14C8
    x"C0",x"90",x"05",x"B9",x"00",x"10",x"B0",x"03", -- 0x14D0
    x"B9",x"00",x"11",x"91",x"B0",x"88",x"D0",x"EF", -- 0x14D8
    x"20",x"F2",x"8F",x"A0",x"D5",x"A9",x"00",x"91", -- 0x14E0
    x"B0",x"60",x"C9",x"08",x"D0",x"15",x"20",x"11", -- 0x14E8
    x"84",x"A4",x"F0",x"84",x"B0",x"A4",x"F1",x"84", -- 0x14F0
    x"B1",x"A4",x"EF",x"C0",x"7F",x"D0",x"4C",x"4C", -- 0x14F8
    x"13",x"B9",x"00",x"4C",x"F6",x"A0",x"00",x"00", -- 0x1500
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1508
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1510
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1518
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1520
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1528
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1530
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1538
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x1540
    x"00",x"00",x"00",x"C0",x"7D",x"90",x"2B",x"20", -- 0x1548
    x"4D",x"83",x"20",x"47",x"83",x"C0",x"7E",x"F0", -- 0x1550
    x"09",x"A0",x"00",x"AD",x"04",x"0F",x"91",x"B0", -- 0x1558
    x"98",x"60",x"A9",x"00",x"A8",x"91",x"B0",x"C8", -- 0x1560
    x"AD",x"07",x"0F",x"91",x"B0",x"C8",x"AD",x"06", -- 0x1568
    x"0F",x"29",x"03",x"91",x"B0",x"C8",x"A9",x"00", -- 0x1570
    x"91",x"B0",x"60",x"20",x"11",x"84",x"48",x"20", -- 0x1578
    x"62",x"82",x"86",x"B0",x"8E",x"DC",x"10",x"84", -- 0x1580
    x"B1",x"8C",x"DD",x"10",x"A2",x"00",x"A0",x"00", -- 0x1588
    x"20",x"EA",x"80",x"20",x"DA",x"80",x"C0",x"12", -- 0x1590
    x"D0",x"F9",x"68",x"AA",x"E8",x"E0",x"08",x"B0", -- 0x1598
    x"08",x"BD",x"8C",x"99",x"48",x"BD",x"84",x"99", -- 0x15A0
    x"48",x"60",x"C9",x"09",x"B0",x"FB",x"86",x"B5", -- 0x15A8
    x"AA",x"BD",x"75",x"99",x"48",x"BD",x"6C",x"99", -- 0x15B0
    x"48",x"8A",x"A6",x"B5",x"60",x"A9",x"FF",x"95", -- 0x15B8
    x"02",x"95",x"03",x"AD",x"DA",x"10",x"95",x"00", -- 0x15C0
    x"AD",x"DB",x"10",x"95",x"01",x"A9",x"00",x"60", -- 0x15C8
    x"C9",x"09",x"B0",x"FB",x"20",x"E1",x"83",x"8E", -- 0x15D0
    x"7D",x"10",x"8C",x"7E",x"10",x"A8",x"BA",x"A9", -- 0x15D8
    x"00",x"4C",x"D8",x"A0",x"B9",x"AB",x"99",x"8D", -- 0x15E0
    x"D8",x"10",x"B9",x"B4",x"99",x"8D",x"D9",x"10", -- 0x15E8
    x"B9",x"BD",x"99",x"4A",x"08",x"4A",x"08",x"8D", -- 0x15F0
    x"7F",x"10",x"20",x"56",x"97",x"A0",x"0C",x"B1", -- 0x15F8
    x"B4",x"99",x"60",x"10",x"88",x"10",x"F8",x"AD", -- 0x1600
    x"63",x"10",x"2D",x"64",x"10",x"0D",x"D7",x"10", -- 0x1608
    x"18",x"69",x"01",x"4C",x"EB",x"A0",x"EA",x"8D", -- 0x1610
    x"81",x"10",x"AD",x"7F",x"10",x"B0",x"07",x"A2", -- 0x1618
    x"61",x"A0",x"10",x"20",x"06",x"04",x"28",x"B0", -- 0x1620
    x"04",x"28",x"6C",x"D8",x"10",x"A2",x"03",x"BD", -- 0x1628
    x"69",x"10",x"95",x"B6",x"CA",x"10",x"F8",x"A2", -- 0x1630
    x"B6",x"AC",x"60",x"10",x"A9",x"00",x"28",x"B0", -- 0x1638
    x"03",x"20",x"A7",x"92",x"20",x"2E",x"90",x"A2", -- 0x1640
    x"03",x"B5",x"B6",x"9D",x"69",x"10",x"CA",x"10", -- 0x1648
    x"F8",x"20",x"48",x"97",x"30",x"0D",x"AC",x"60", -- 0x1650
    x"10",x"20",x"2A",x"96",x"B0",x"0D",x"A2",x"09", -- 0x1658
    x"20",x"3C",x"97",x"A2",x"05",x"20",x"3C",x"97", -- 0x1660
    x"D0",x"EC",x"18",x"08",x"20",x"48",x"97",x"A2", -- 0x1668
    x"05",x"20",x"3C",x"97",x"A0",x"0C",x"20",x"56", -- 0x1670
    x"97",x"B9",x"60",x"10",x"91",x"B4",x"88",x"10", -- 0x1678
    x"F8",x"28",x"60",x"20",x"4D",x"83",x"20",x"4D", -- 0x1680
    x"AB",x"A9",x"95",x"8D",x"D8",x"10",x"A9",x"96", -- 0x1688
    x"8D",x"D9",x"10",x"D0",x"BC",x"AC",x"69",x"10", -- 0x1690
    x"CC",x"05",x"0F",x"B0",x"28",x"B9",x"0F",x"0E", -- 0x1698
    x"20",x"EE",x"82",x"45",x"CE",x"B0",x"02",x"29", -- 0x16A0
    x"DF",x"29",x"7F",x"F0",x"05",x"20",x"10",x"82", -- 0x16A8
    x"D0",x"E6",x"A9",x"07",x"20",x"6A",x"97",x"85", -- 0x16B0
    x"B0",x"B9",x"08",x"0E",x"20",x"6A",x"97",x"C8", -- 0x16B8
    x"C6",x"B0",x"D0",x"F5",x"18",x"8C",x"69",x"10", -- 0x16C0
    x"AD",x"04",x"0F",x"8D",x"60",x"10",x"60",x"20", -- 0x16C8
    x"4D",x"83",x"20",x"4D",x"AB",x"A9",x"0C",x"20", -- 0x16D0
    x"6A",x"97",x"A0",x"00",x"B9",x"00",x"0E",x"20", -- 0x16D8
    x"6A",x"97",x"C8",x"C0",x"08",x"D0",x"F5",x"B9", -- 0x16E0
    x"F8",x"0E",x"20",x"6A",x"97",x"C8",x"C0",x"0C", -- 0x16E8
    x"D0",x"F5",x"AD",x"06",x"0F",x"20",x"05",x"82", -- 0x16F0
    x"20",x"6A",x"97",x"A5",x"CF",x"4C",x"6A",x"97", -- 0x16F8
    x"20",x"61",x"97",x"AD",x"CB",x"10",x"09",x"30", -- 0x1700
    x"20",x"6A",x"97",x"20",x"61",x"97",x"AD",x"CA", -- 0x1708
    x"10",x"4C",x"6A",x"97",x"20",x"61",x"97",x"AD", -- 0x1710
    x"CD",x"10",x"09",x"30",x"20",x"6A",x"97",x"20", -- 0x1718
    x"61",x"97",x"AD",x"CC",x"10",x"4C",x"6A",x"97", -- 0x1720
    x"48",x"AD",x"61",x"10",x"85",x"B8",x"AD",x"62", -- 0x1728
    x"10",x"85",x"B9",x"A2",x"00",x"68",x"60",x"20", -- 0x1730
    x"E1",x"83",x"A2",x"01",x"A0",x"04",x"FE",x"60", -- 0x1738
    x"10",x"D0",x"04",x"E8",x"88",x"D0",x"F7",x"60", -- 0x1740
    x"A2",x"03",x"A9",x"FF",x"5D",x"65",x"10",x"9D", -- 0x1748
    x"65",x"10",x"CA",x"10",x"F5",x"60",x"AD",x"7D", -- 0x1750
    x"10",x"85",x"B4",x"AD",x"7E",x"10",x"85",x"B5", -- 0x1758
    x"60",x"A9",x"01",x"D0",x"05",x"20",x"C1",x"90", -- 0x1760
    x"B0",x"F6",x"2C",x"81",x"10",x"10",x"06",x"8D", -- 0x1768
    x"E5",x"FE",x"4C",x"37",x"97",x"20",x"28",x"97", -- 0x1770
    x"81",x"B8",x"4C",x"37",x"97",x"20",x"85",x"97", -- 0x1778
    x"20",x"AA",x"91",x"18",x"60",x"2C",x"81",x"10", -- 0x1780
    x"10",x"06",x"AD",x"E5",x"FE",x"4C",x"37",x"97", -- 0x1788
    x"20",x"28",x"97",x"A1",x"B8",x"4C",x"37",x"97", -- 0x1790
    x"2C",x"C8",x"10",x"30",x"03",x"CE",x"C8",x"10", -- 0x1798
    x"60",x"20",x"5A",x"98",x"20",x"7E",x"83",x"A9", -- 0x17A0
    x"01",x"60",x"20",x"37",x"98",x"20",x"7E",x"83", -- 0x17A8
    x"20",x"D1",x"82",x"90",x"24",x"20",x"37",x"98", -- 0x17B0
    x"20",x"DF",x"97",x"20",x"FB",x"97",x"50",x"16", -- 0x17B8
    x"20",x"37",x"98",x"20",x"DF",x"97",x"50",x"11", -- 0x17C0
    x"20",x"37",x"98",x"20",x"FB",x"97",x"50",x"09", -- 0x17C8
    x"20",x"5A",x"98",x"20",x"4F",x"98",x"20",x"1E", -- 0x17D0
    x"98",x"20",x"C3",x"88",x"A9",x"01",x"60",x"20", -- 0x17D8
    x"E1",x"83",x"A0",x"02",x"B1",x"B0",x"9D",x"08", -- 0x17E0
    x"0F",x"C8",x"B1",x"B0",x"9D",x"09",x"0F",x"C8", -- 0x17E8
    x"B1",x"B0",x"0A",x"0A",x"5D",x"0E",x"0F",x"29", -- 0x17F0
    x"0C",x"10",x"1B",x"20",x"E1",x"83",x"A0",x"06", -- 0x17F8
    x"B1",x"B0",x"9D",x"0A",x"0F",x"C8",x"B1",x"B0", -- 0x1800
    x"9D",x"0B",x"0F",x"C8",x"B1",x"B0",x"6A",x"6A", -- 0x1808
    x"6A",x"5D",x"0E",x"0F",x"29",x"C0",x"5D",x"0E", -- 0x1810
    x"0F",x"9D",x"0E",x"0F",x"B8",x"60",x"20",x"E1", -- 0x1818
    x"83",x"A0",x"0E",x"B1",x"B0",x"29",x"0A",x"F0", -- 0x1820
    x"02",x"A9",x"80",x"5D",x"0F",x"0E",x"29",x"80", -- 0x1828
    x"5D",x"0F",x"0E",x"9D",x"0F",x"0E",x"60",x"20", -- 0x1830
    x"64",x"98",x"90",x"23",x"B9",x"0F",x"0E",x"10", -- 0x1838
    x"22",x"20",x"2B",x"80",x"C3",x"6C",x"6F",x"63", -- 0x1840
    x"6B",x"65",x"64",x"00",x"20",x"3C",x"98",x"20", -- 0x1848
    x"E1",x"83",x"20",x"9E",x"8F",x"90",x"21",x"4C", -- 0x1850
    x"02",x"8F",x"20",x"64",x"98",x"B0",x"19",x"68", -- 0x1858
    x"68",x"A9",x"00",x"60",x"20",x"06",x"81",x"20", -- 0x1860
    x"96",x"82",x"90",x"0C",x"98",x"AA",x"AD",x"DC", -- 0x1868
    x"10",x"85",x"B0",x"AD",x"DD",x"10",x"85",x"B1", -- 0x1870
    x"60",x"A9",x"83",x"20",x"F4",x"FF",x"8C",x"D0", -- 0x1878
    x"10",x"A9",x"84",x"20",x"F4",x"FF",x"98",x"38", -- 0x1880
    x"ED",x"D0",x"10",x"8D",x"D1",x"10",x"60",x"A2", -- 0x1888
    x"0A",x"20",x"2C",x"99",x"20",x"9E",x"98",x"A0", -- 0x1890
    x"D5",x"A9",x"FF",x"91",x"B0",x"60",x"48",x"A6", -- 0x1898
    x"F4",x"A9",x"00",x"85",x"B0",x"BD",x"F0",x"0D", -- 0x18A0
    x"85",x"B1",x"68",x"60",x"00",x"00",x"00",x"00", -- 0x18A8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18B0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18B8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18C0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18C8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18D0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18D8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18E0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18E8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x18F8
    x"00",x"00",x"00",x"00",x"00",x"60",x"20",x"E1", -- 0x1900
    x"83",x"A9",x"0F",x"A2",x"01",x"A0",x"00",x"F0", -- 0x1908
    x"25",x"A9",x"C7",x"A2",x"00",x"F0",x"F6",x"AA", -- 0x1910
    x"A9",x"03",x"D0",x"1A",x"A9",x"EC",x"D0",x"12", -- 0x1918
    x"A9",x"C7",x"D0",x"0E",x"A9",x"EA",x"D0",x"0A", -- 0x1920
    x"A9",x"A8",x"D0",x"06",x"A9",x"8F",x"D0",x"06", -- 0x1928
    x"A9",x"FF",x"A2",x"00",x"A0",x"FF",x"4C",x"F4", -- 0x1930
    x"FF",x"4C",x"2E",x"21",x"42",x"4F",x"4F",x"54", -- 0x1938
    x"0D",x"45",x"2E",x"21",x"42",x"4F",x"4F",x"54", -- 0x1940
    x"0D",x"1B",x"FF",x"1E",x"FF",x"21",x"FF",x"24", -- 0x1948
    x"FF",x"27",x"FF",x"2A",x"FF",x"2D",x"FF",x"7B", -- 0x1950
    x"95",x"00",x"07",x"90",x"00",x"C1",x"90",x"00", -- 0x1958
    x"AA",x"91",x"00",x"D0",x"95",x"00",x"93",x"8E", -- 0x1960
    x"00",x"AA",x"95",x"00",x"1B",x"8C",x"D3",x"6B", -- 0x1968
    x"D3",x"1D",x"E1",x"DC",x"97",x"89",x"90",x"87", -- 0x1970
    x"86",x"87",x"84",x"8D",x"8D",x"97",x"F1",x"3C", -- 0x1978
    x"BC",x"8F",x"9B",x"95",x"93",x"85",x"B4",x"BF", -- 0x1980
    x"C7",x"CF",x"A0",x"A9",x"87",x"87",x"97",x"97", -- 0x1988
    x"97",x"97",x"97",x"97",x"12",x"32",x"5D",x"CD", -- 0x1990
    x"A2",x"BD",x"87",x"8D",x"8D",x"8D",x"8D",x"8D", -- 0x1998
    x"8D",x"8D",x"74",x"54",x"00",x"0F",x"1A",x"0F", -- 0x19A0
    x"1A",x"63",x"43",x"B7",x"7D",x"7D",x"65",x"65", -- 0x19A8
    x"CF",x"00",x"14",x"83",x"85",x"97",x"97",x"97", -- 0x19B0
    x"97",x"96",x"97",x"97",x"96",x"04",x"02",x"03", -- 0x19B8
    x"06",x"07",x"04",x"04",x"04",x"04",x"98",x"A2", -- 0x19C0
    x"FF",x"A0",x"0E",x"48",x"20",x"65",x"80",x"0D", -- 0x19C8
    x"44",x"46",x"53",x"20",x"30",x"2E",x"39",x"30", -- 0x19D0
    x"0D",x"86",x"B8",x"20",x"CB",x"9F",x"20",x"19", -- 0x19D8
    x"9A",x"20",x"9A",x"9F",x"88",x"D0",x"F4",x"68", -- 0x19E0
    x"A8",x"A2",x"A0",x"4C",x"71",x"86",x"98",x"A2", -- 0x19E8
    x"74",x"A0",x"05",x"D0",x"D6",x"20",x"BF",x"86", -- 0x19F0
    x"F0",x"60",x"20",x"C5",x"FF",x"90",x"FB",x"B0", -- 0x19F8
    x"E8",x"20",x"BF",x"86",x"D0",x"54",x"20",x"33", -- 0x1A00
    x"80",x"DC",x"53",x"79",x"6E",x"74",x"61",x"78", -- 0x1A08
    x"3A",x"20",x"EA",x"20",x"19",x"9A",x"4C",x"8A", -- 0x1A10
    x"80",x"A6",x"B8",x"E8",x"BD",x"B8",x"85",x"30", -- 0x1A18
    x"06",x"20",x"9C",x"80",x"4C",x"1B",x"9A",x"E8", -- 0x1A20
    x"E8",x"86",x"B8",x"BD",x"B8",x"85",x"20",x"34", -- 0x1A28
    x"9A",x"20",x"05",x"82",x"20",x"E1",x"83",x"29", -- 0x1A30
    x"0F",x"F0",x"1F",x"A8",x"A9",x"20",x"20",x"9C", -- 0x1A38
    x"80",x"A2",x"00",x"BD",x"5B",x"9A",x"F0",x"03", -- 0x1A40
    x"E8",x"D0",x"F8",x"88",x"D0",x"FA",x"E8",x"BD", -- 0x1A48
    x"5B",x"9A",x"F0",x"06",x"20",x"9C",x"80",x"4C", -- 0x1A50
    x"4E",x"9A",x"60",x"00",x"3C",x"66",x"73",x"70", -- 0x1A58
    x"3E",x"00",x"3C",x"61",x"66",x"73",x"70",x"3E", -- 0x1A60
    x"00",x"28",x"4C",x"29",x"00",x"3C",x"73",x"72", -- 0x1A68
    x"63",x"20",x"64",x"72",x"76",x"3E",x"00",x"3C", -- 0x1A70
    x"64",x"65",x"73",x"74",x"20",x"64",x"72",x"76", -- 0x1A78
    x"3E",x"00",x"3C",x"64",x"65",x"73",x"74",x"20", -- 0x1A80
    x"64",x"72",x"76",x"3E",x"20",x"3C",x"61",x"66", -- 0x1A88
    x"73",x"70",x"3E",x"00",x"3C",x"6F",x"6C",x"64", -- 0x1A90
    x"20",x"66",x"73",x"70",x"3E",x"00",x"3C",x"6E", -- 0x1A98
    x"65",x"77",x"20",x"66",x"73",x"70",x"3E",x"00", -- 0x1AA0
    x"28",x"3C",x"64",x"69",x"72",x"3E",x"29",x"00", -- 0x1AA8
    x"28",x"3C",x"64",x"72",x"76",x"3E",x"29",x"00", -- 0x1AB0
    x"3C",x"74",x"69",x"74",x"6C",x"65",x"3E",x"00", -- 0x1AB8
    x"20",x"58",x"83",x"20",x"65",x"80",x"43",x"6F", -- 0x1AC0
    x"6D",x"70",x"61",x"63",x"74",x"69",x"6E",x"67", -- 0x1AC8
    x"20",x"64",x"72",x"69",x"76",x"65",x"20",x"8D", -- 0x1AD0
    x"D2",x"10",x"8D",x"D3",x"10",x"20",x"CA",x"80", -- 0x1AD8
    x"20",x"9A",x"9F",x"A0",x"00",x"20",x"05",x"8E", -- 0x1AE0
    x"20",x"79",x"98",x"20",x"47",x"83",x"AC",x"05", -- 0x1AE8
    x"0F",x"84",x"CC",x"A9",x"02",x"85",x"CA",x"A9", -- 0x1AF0
    x"00",x"85",x"CB",x"A4",x"CC",x"20",x"19",x"82", -- 0x1AF8
    x"C0",x"F8",x"D0",x"3C",x"20",x"65",x"80",x"44", -- 0x1B00
    x"69",x"73",x"6B",x"20",x"63",x"6F",x"6D",x"70", -- 0x1B08
    x"61",x"63",x"74",x"65",x"64",x"20",x"EA",x"38", -- 0x1B10
    x"AD",x"07",x"0F",x"E5",x"CA",x"48",x"AD",x"06", -- 0x1B18
    x"0F",x"29",x"03",x"E5",x"CB",x"20",x"CA",x"80", -- 0x1B20
    x"68",x"20",x"C2",x"80",x"20",x"65",x"80",x"20", -- 0x1B28
    x"66",x"72",x"65",x"65",x"20",x"73",x"65",x"63", -- 0x1B30
    x"74",x"6F",x"72",x"73",x"0D",x"A9",x"04",x"60", -- 0x1B38
    x"84",x"CC",x"20",x"FC",x"82",x"A4",x"CC",x"B9", -- 0x1B40
    x"0E",x"0F",x"29",x"30",x"19",x"0D",x"0F",x"19", -- 0x1B48
    x"0C",x"0F",x"F0",x"61",x"A9",x"00",x"85",x"BE", -- 0x1B50
    x"85",x"C2",x"A9",x"FF",x"18",x"79",x"0C",x"0F", -- 0x1B58
    x"A9",x"00",x"79",x"0D",x"0F",x"85",x"C6",x"B9", -- 0x1B60
    x"0E",x"0F",x"08",x"20",x"FD",x"81",x"28",x"69", -- 0x1B68
    x"00",x"85",x"C7",x"B9",x"0F",x"0F",x"85",x"C8", -- 0x1B70
    x"B9",x"0E",x"0F",x"29",x"03",x"85",x"C9",x"C5", -- 0x1B78
    x"CB",x"D0",x"14",x"A5",x"C8",x"C5",x"CA",x"D0", -- 0x1B80
    x"0E",x"18",x"65",x"C6",x"85",x"CA",x"A5",x"CB", -- 0x1B88
    x"65",x"C7",x"85",x"CB",x"4C",x"B5",x"9B",x"A5", -- 0x1B90
    x"CA",x"99",x"0F",x"0F",x"B9",x"0E",x"0F",x"29", -- 0x1B98
    x"FC",x"05",x"CB",x"99",x"0E",x"0F",x"A9",x"00", -- 0x1BA0
    x"85",x"A8",x"85",x"A9",x"20",x"B4",x"8A",x"20", -- 0x1BA8
    x"06",x"9E",x"20",x"47",x"83",x"A4",x"CC",x"20", -- 0x1BB0
    x"01",x"83",x"4C",x"FB",x"9A",x"2C",x"C8",x"10", -- 0x1BB8
    x"10",x"75",x"20",x"33",x"80",x"BD",x"4E",x"6F", -- 0x1BC0
    x"74",x"20",x"65",x"6E",x"61",x"62",x"6C",x"65", -- 0x1BC8
    x"64",x"00",x"20",x"BF",x"86",x"D0",x"03",x"4C", -- 0x1BD0
    x"06",x"9A",x"20",x"5D",x"83",x"8D",x"D2",x"10", -- 0x1BD8
    x"20",x"BF",x"86",x"F0",x"F2",x"20",x"5D",x"83", -- 0x1BE0
    x"8D",x"D3",x"10",x"98",x"48",x"A9",x"00",x"85", -- 0x1BE8
    x"A9",x"AD",x"D3",x"10",x"CD",x"D2",x"10",x"D0", -- 0x1BF0
    x"06",x"A9",x"FF",x"85",x"A9",x"85",x"AA",x"20", -- 0x1BF8
    x"79",x"98",x"20",x"65",x"80",x"43",x"6F",x"70", -- 0x1C00
    x"79",x"69",x"6E",x"67",x"20",x"66",x"72",x"6F", -- 0x1C08
    x"6D",x"20",x"64",x"72",x"69",x"76",x"65",x"20", -- 0x1C10
    x"AD",x"D2",x"10",x"20",x"CA",x"80",x"20",x"65", -- 0x1C18
    x"80",x"20",x"74",x"6F",x"20",x"64",x"72",x"69", -- 0x1C20
    x"76",x"65",x"20",x"AD",x"D3",x"10",x"20",x"CA", -- 0x1C28
    x"80",x"20",x"9A",x"9F",x"68",x"A8",x"18",x"60", -- 0x1C30
    x"20",x"E1",x"83",x"24",x"A9",x"10",x"0B",x"A9", -- 0x1C38
    x"00",x"F0",x"0A",x"20",x"E1",x"83",x"24",x"A9", -- 0x1C40
    x"30",x"01",x"60",x"A9",x"80",x"C5",x"AA",x"F0", -- 0x1C48
    x"F9",x"85",x"AA",x"20",x"65",x"80",x"49",x"6E", -- 0x1C50
    x"73",x"65",x"72",x"74",x"20",x"EA",x"24",x"AA", -- 0x1C58
    x"30",x"0B",x"20",x"65",x"80",x"73",x"6F",x"75", -- 0x1C60
    x"72",x"63",x"65",x"90",x"0F",x"20",x"65",x"80", -- 0x1C68
    x"64",x"65",x"73",x"74",x"69",x"6E",x"61",x"74", -- 0x1C70
    x"69",x"6F",x"6E",x"EA",x"20",x"65",x"80",x"20", -- 0x1C78
    x"64",x"69",x"73",x"6B",x"20",x"61",x"6E",x"64", -- 0x1C80
    x"20",x"68",x"69",x"74",x"20",x"61",x"20",x"6B", -- 0x1C88
    x"65",x"79",x"EA",x"20",x"06",x"99",x"20",x"E0", -- 0x1C90
    x"FF",x"B0",x"19",x"4C",x"9A",x"9F",x"20",x"06", -- 0x1C98
    x"99",x"20",x"E0",x"FF",x"B0",x"0E",x"29",x"5F", -- 0x1CA0
    x"C9",x"59",x"08",x"F0",x"02",x"A9",x"4E",x"20", -- 0x1CA8
    x"9C",x"80",x"28",x"60",x"A6",x"B6",x"9A",x"60", -- 0x1CB0
    x"4C",x"58",x"89",x"20",x"BD",x"9B",x"20",x"D2", -- 0x1CB8
    x"9B",x"A9",x"00",x"85",x"C9",x"85",x"CB",x"85", -- 0x1CC0
    x"CA",x"85",x"C8",x"85",x"A8",x"20",x"38",x"9C", -- 0x1CC8
    x"AD",x"D2",x"10",x"85",x"CF",x"20",x"4D",x"AB", -- 0x1CD0
    x"AD",x"07",x"0F",x"85",x"C6",x"AD",x"06",x"0F", -- 0x1CD8
    x"29",x"03",x"85",x"C7",x"AD",x"06",x"0F",x"29", -- 0x1CE0
    x"F0",x"8D",x"D8",x"10",x"20",x"43",x"9C",x"AD", -- 0x1CE8
    x"D3",x"10",x"85",x"CF",x"20",x"4D",x"AB",x"AD", -- 0x1CF0
    x"06",x"0F",x"29",x"03",x"C5",x"C7",x"90",x"B8", -- 0x1CF8
    x"D0",x"07",x"AD",x"07",x"0F",x"C5",x"C6",x"90", -- 0x1D00
    x"AF",x"20",x"06",x"9E",x"AD",x"06",x"0F",x"48", -- 0x1D08
    x"AD",x"07",x"0F",x"48",x"20",x"4D",x"AB",x"68", -- 0x1D10
    x"8D",x"07",x"0F",x"68",x"29",x"0F",x"0D",x"D8", -- 0x1D18
    x"10",x"8D",x"06",x"0F",x"4C",x"B4",x"8A",x"20", -- 0x1D20
    x"5E",x"82",x"20",x"D2",x"9B",x"20",x"BF",x"86", -- 0x1D28
    x"D0",x"03",x"4C",x"06",x"9A",x"20",x"FE",x"80", -- 0x1D30
    x"20",x"38",x"9C",x"AD",x"D2",x"10",x"20",x"7E", -- 0x1D38
    x"87",x"20",x"96",x"82",x"B0",x"03",x"4C",x"76", -- 0x1D40
    x"82",x"84",x"AB",x"20",x"01",x"83",x"A2",x"00", -- 0x1D48
    x"B5",x"C7",x"9D",x"58",x"10",x"B9",x"08",x"0E", -- 0x1D50
    x"95",x"C7",x"9D",x"50",x"10",x"B9",x"08",x"0F", -- 0x1D58
    x"95",x"BD",x"9D",x"47",x"10",x"E8",x"C8",x"E0", -- 0x1D60
    x"08",x"D0",x"E5",x"A5",x"C3",x"20",x"FD",x"81", -- 0x1D68
    x"85",x"C5",x"A5",x"C1",x"18",x"69",x"FF",x"A5", -- 0x1D70
    x"C2",x"69",x"00",x"85",x"C6",x"A5",x"C5",x"69", -- 0x1D78
    x"00",x"85",x"C7",x"AD",x"4E",x"10",x"85",x"C8", -- 0x1D80
    x"AD",x"4D",x"10",x"29",x"03",x"85",x"C9",x"A9", -- 0x1D88
    x"FF",x"85",x"A8",x"20",x"06",x"9E",x"20",x"38", -- 0x1D90
    x"9C",x"AD",x"D2",x"10",x"20",x"7E",x"87",x"20", -- 0x1D98
    x"47",x"83",x"A2",x"07",x"BD",x"58",x"10",x"95", -- 0x1DA0
    x"C7",x"CA",x"10",x"F8",x"A4",x"AB",x"8C",x"CE", -- 0x1DA8
    x"10",x"20",x"9D",x"82",x"B0",x"93",x"60",x"20", -- 0x1DB0
    x"F5",x"9D",x"20",x"43",x"9C",x"AD",x"D3",x"10", -- 0x1DB8
    x"85",x"CF",x"A5",x"CE",x"48",x"20",x"47",x"83", -- 0x1DC0
    x"20",x"96",x"82",x"90",x"03",x"20",x"D1",x"82", -- 0x1DC8
    x"68",x"85",x"CE",x"20",x"3F",x"8A",x"20",x"56", -- 0x1DD0
    x"8A",x"A5",x"C4",x"20",x"FD",x"81",x"85",x"C6", -- 0x1DD8
    x"20",x"9D",x"89",x"A5",x"C4",x"29",x"03",x"48", -- 0x1DE0
    x"A5",x"C5",x"48",x"20",x"F5",x"9D",x"68",x"85", -- 0x1DE8
    x"CA",x"68",x"85",x"CB",x"60",x"A2",x"11",x"BD", -- 0x1DF0
    x"45",x"10",x"B4",x"BC",x"95",x"BC",x"98",x"9D", -- 0x1DF8
    x"45",x"10",x"CA",x"10",x"F2",x"60",x"20",x"8D", -- 0x1E00
    x"A0",x"A9",x"00",x"85",x"BE",x"85",x"C2",x"A5", -- 0x1E08
    x"C6",x"A8",x"CD",x"D1",x"10",x"A5",x"C7",x"E9", -- 0x1E10
    x"00",x"90",x"03",x"AC",x"D1",x"10",x"84",x"C3", -- 0x1E18
    x"A5",x"C8",x"85",x"C5",x"A5",x"C9",x"85",x"C4", -- 0x1E20
    x"AD",x"D0",x"10",x"85",x"BF",x"AD",x"D2",x"10", -- 0x1E28
    x"85",x"CF",x"20",x"38",x"9C",x"20",x"0B",x"B9", -- 0x1E30
    x"20",x"C6",x"87",x"AD",x"D3",x"10",x"85",x"CF", -- 0x1E38
    x"24",x"A8",x"10",x"07",x"20",x"B7",x"9D",x"A9", -- 0x1E40
    x"00",x"85",x"A8",x"A5",x"CA",x"85",x"C5",x"A5", -- 0x1E48
    x"CB",x"85",x"C4",x"AD",x"D0",x"10",x"85",x"BF", -- 0x1E50
    x"20",x"43",x"9C",x"20",x"0B",x"B9",x"20",x"8F", -- 0x1E58
    x"87",x"A5",x"C3",x"18",x"65",x"CA",x"85",x"CA", -- 0x1E60
    x"90",x"02",x"E6",x"CB",x"A5",x"C3",x"18",x"65", -- 0x1E68
    x"C8",x"85",x"C8",x"90",x"02",x"E6",x"C9",x"38", -- 0x1E70
    x"A5",x"C6",x"E5",x"C3",x"85",x"C6",x"B0",x"02", -- 0x1E78
    x"C6",x"C7",x"05",x"C7",x"D0",x"89",x"60",x"20", -- 0x1E80
    x"D7",x"9F",x"A9",x"00",x"F0",x"05",x"20",x"D7", -- 0x1E88
    x"9F",x"A9",x"FF",x"85",x"AB",x"A9",x"C0",x"20", -- 0x1E90
    x"CE",x"FF",x"A8",x"A9",x"0D",x"C0",x"00",x"D0", -- 0x1E98
    x"1E",x"4C",x"76",x"82",x"20",x"D7",x"FF",x"B0", -- 0x1EA0
    x"1E",x"C9",x"0A",x"F0",x"F7",x"28",x"D0",x"08", -- 0x1EA8
    x"48",x"20",x"A2",x"9F",x"20",x"CE",x"9F",x"68", -- 0x1EB0
    x"20",x"E3",x"FF",x"24",x"FF",x"30",x"09",x"25", -- 0x1EB8
    x"AB",x"C9",x"0D",x"08",x"4C",x"A4",x"9E",x"28", -- 0x1EC0
    x"20",x"9A",x"9F",x"A9",x"00",x"4C",x"CE",x"FF", -- 0x1EC8
    x"20",x"D7",x"9F",x"A9",x"C0",x"20",x"CE",x"FF", -- 0x1ED0
    x"A8",x"F0",x"C6",x"A6",x"F4",x"BD",x"F0",x"0D", -- 0x1ED8
    x"85",x"AD",x"E6",x"AD",x"24",x"FF",x"30",x"E3", -- 0x1EE0
    x"A5",x"A9",x"20",x"C2",x"80",x"A5",x"A8",x"20", -- 0x1EE8
    x"C2",x"80",x"20",x"CE",x"9F",x"A9",x"07",x"85", -- 0x1EF0
    x"AC",x"A2",x"00",x"20",x"D7",x"FF",x"B0",x"0D", -- 0x1EF8
    x"81",x"AC",x"20",x"C2",x"80",x"20",x"CE",x"9F", -- 0x1F00
    x"C6",x"AC",x"10",x"EF",x"18",x"08",x"90",x"0E", -- 0x1F08
    x"20",x"65",x"80",x"2A",x"2A",x"20",x"A9",x"00", -- 0x1F10
    x"81",x"AC",x"C6",x"AC",x"10",x"F2",x"A9",x"07", -- 0x1F18
    x"85",x"AC",x"A1",x"AC",x"C9",x"7F",x"B0",x"04", -- 0x1F20
    x"C9",x"20",x"B0",x"02",x"A9",x"2E",x"20",x"E3", -- 0x1F28
    x"FF",x"C6",x"AC",x"10",x"ED",x"20",x"9A",x"9F", -- 0x1F30
    x"A9",x"08",x"18",x"65",x"A8",x"85",x"A8",x"90", -- 0x1F38
    x"02",x"E6",x"A9",x"28",x"90",x"9E",x"B0",x"83", -- 0x1F40
    x"20",x"D7",x"9F",x"A9",x"80",x"20",x"CE",x"FF", -- 0x1F48
    x"85",x"AB",x"20",x"A2",x"9F",x"20",x"CE",x"9F", -- 0x1F50
    x"A6",x"F4",x"BC",x"F0",x"0D",x"C8",x"84",x"AD", -- 0x1F58
    x"A2",x"AC",x"A0",x"FF",x"84",x"AE",x"84",x"B0", -- 0x1F60
    x"C8",x"84",x"AC",x"84",x"AF",x"98",x"20",x"F1", -- 0x1F68
    x"FF",x"08",x"84",x"AA",x"A4",x"AB",x"A2",x"00", -- 0x1F70
    x"F0",x"07",x"A1",x"AC",x"20",x"D4",x"FF",x"E6", -- 0x1F78
    x"AC",x"A5",x"AC",x"C5",x"AA",x"D0",x"F3",x"28", -- 0x1F80
    x"B0",x"08",x"A9",x"0D",x"20",x"D4",x"FF",x"4C", -- 0x1F88
    x"52",x"9F",x"A9",x"7E",x"20",x"F4",x"FF",x"20", -- 0x1F90
    x"CB",x"9E",x"48",x"A9",x"0D",x"20",x"9C",x"80", -- 0x1F98
    x"68",x"60",x"F8",x"18",x"A5",x"A8",x"69",x"01", -- 0x1FA0
    x"85",x"A8",x"A5",x"A9",x"69",x"00",x"85",x"A9", -- 0x1FA8
    x"D8",x"18",x"20",x"B7",x"9F",x"A5",x"A8",x"48", -- 0x1FB0
    x"08",x"20",x"05",x"82",x"28",x"20",x"C1",x"9F", -- 0x1FB8
    x"68",x"AA",x"B0",x"02",x"F0",x"08",x"20",x"CA", -- 0x1FC0
    x"80",x"38",x"60",x"20",x"CE",x"9F",x"48",x"A9", -- 0x1FC8
    x"20",x"20",x"9C",x"80",x"68",x"18",x"60",x"BA", -- 0x1FD0
    x"A9",x"00",x"9D",x"07",x"01",x"88",x"C8",x"B1", -- 0x1FD8
    x"F2",x"C9",x"20",x"F0",x"F9",x"C9",x"0D",x"D0", -- 0x1FE0
    x"03",x"4C",x"06",x"9A",x"A9",x"00",x"85",x"A8", -- 0x1FE8
    x"85",x"A9",x"48",x"98",x"18",x"65",x"F2",x"AA", -- 0x1FF0
    x"A5",x"F3",x"69",x"00",x"A8",x"68",x"60",x"6D", -- 0x1FF8
    x"20",x"7B",x"A1",x"68",x"85",x"B8",x"68",x"85", -- 0x2000
    x"B9",x"20",x"0F",x"A0",x"4C",x"00",x"01",x"A0", -- 0x2008
    x"00",x"8C",x"00",x"01",x"C8",x"F0",x"07",x"B1", -- 0x2010
    x"B8",x"99",x"00",x"01",x"D0",x"F6",x"60",x"A2", -- 0x2018
    x"FF",x"D0",x"02",x"A2",x"00",x"A0",x"FF",x"8C", -- 0x2020
    x"82",x"10",x"85",x"B0",x"86",x"B1",x"8D",x"02", -- 0x2028
    x"0D",x"20",x"7B",x"A1",x"68",x"85",x"B8",x"68", -- 0x2030
    x"85",x"B9",x"20",x"0F",x"A0",x"A5",x"B0",x"20", -- 0x2038
    x"69",x"A0",x"A5",x"B1",x"F0",x"1B",x"A9",x"2F", -- 0x2040
    x"99",x"00",x"01",x"C8",x"AE",x"41",x"0D",x"BD", -- 0x2048
    x"44",x"0D",x"20",x"69",x"A0",x"BD",x"45",x"0D", -- 0x2050
    x"20",x"69",x"A0",x"BD",x"46",x"0D",x"20",x"69", -- 0x2058
    x"A0",x"A9",x"00",x"99",x"00",x"01",x"4C",x"00", -- 0x2060
    x"01",x"48",x"4A",x"4A",x"4A",x"4A",x"20",x"74", -- 0x2068
    x"A0",x"68",x"29",x"0F",x"18",x"69",x"30",x"C9", -- 0x2070
    x"3A",x"90",x"02",x"69",x"06",x"99",x"00",x"01", -- 0x2078
    x"C8",x"60",x"20",x"00",x"A0",x"11",x"45",x"73", -- 0x2080
    x"63",x"61",x"70",x"65",x"00",x"48",x"A9",x"FF", -- 0x2088
    x"8D",x"74",x"10",x"8D",x"75",x"10",x"68",x"60", -- 0x2090
    x"48",x"A5",x"BE",x"8D",x"72",x"10",x"A5",x"BF", -- 0x2098
    x"8D",x"73",x"10",x"AD",x"74",x"10",x"2D",x"75", -- 0x20A0
    x"10",x"0D",x"D7",x"10",x"49",x"FF",x"8D",x"D6", -- 0x20A8
    x"10",x"38",x"F0",x"0D",x"20",x"C3",x"A0",x"A2", -- 0x20B0
    x"72",x"A0",x"10",x"68",x"48",x"20",x"06",x"04", -- 0x20B8
    x"18",x"68",x"60",x"48",x"A9",x"C1",x"20",x"06", -- 0x20C0
    x"04",x"90",x"F9",x"68",x"60",x"AD",x"D6",x"10", -- 0x20C8
    x"F0",x"05",x"A9",x"81",x"20",x"06",x"04",x"60", -- 0x20D0
    x"9D",x"05",x"01",x"20",x"E4",x"95",x"08",x"AD", -- 0x20D8
    x"81",x"10",x"F0",x"05",x"A9",x"81",x"20",x"06", -- 0x20E0
    x"04",x"28",x"60",x"F0",x"06",x"20",x"C3",x"A0", -- 0x20E8
    x"18",x"A9",x"FF",x"4C",x"17",x"96",x"C9",x"FE", -- 0x20F0
    x"90",x"5A",x"D0",x"1B",x"C0",x"00",x"F0",x"54", -- 0x20F8
    x"A2",x"06",x"A9",x"14",x"20",x"F4",x"FF",x"2C", -- 0x2100
    x"E0",x"FE",x"10",x"FB",x"AD",x"E1",x"FE",x"F0", -- 0x2108
    x"41",x"20",x"EE",x"FF",x"4C",x"07",x"A1",x"A9", -- 0x2110
    x"AD",x"8D",x"20",x"02",x"A9",x"06",x"8D",x"21", -- 0x2118
    x"02",x"A9",x"16",x"8D",x"02",x"02",x"A0",x"00", -- 0x2120
    x"8C",x"03",x"02",x"A9",x"8E",x"8D",x"E0",x"FE", -- 0x2128
    x"B9",x"03",x"8B",x"99",x"00",x"04",x"B9",x"03", -- 0x2130
    x"8C",x"99",x"00",x"05",x"B9",x"03",x"8D",x"99", -- 0x2138
    x"00",x"06",x"88",x"D0",x"EB",x"20",x"21",x"04", -- 0x2140
    x"A2",x"40",x"BD",x"C2",x"8A",x"95",x"16",x"CA", -- 0x2148
    x"10",x"F8",x"A9",x"00",x"60",x"A9",x"FF",x"8D", -- 0x2150
    x"52",x"0D",x"48",x"4C",x"3B",x"93",x"B9",x"14", -- 0x2158
    x"11",x"99",x"10",x"11",x"B9",x"15",x"11",x"99", -- 0x2160
    x"11",x"11",x"B9",x"16",x"11",x"99",x"12",x"11", -- 0x2168
    x"60",x"A2",x"06",x"8E",x"40",x"FE",x"E8",x"8E", -- 0x2170
    x"40",x"FE",x"60",x"A9",x"76",x"4C",x"F4",x"FF", -- 0x2178
    x"A2",x"01",x"A9",x"03",x"8E",x"60",x"FE",x"8D", -- 0x2180
    x"60",x"FE",x"8E",x"60",x"FE",x"8D",x"60",x"FE", -- 0x2188
    x"8E",x"60",x"FE",x"8D",x"60",x"FE",x"8E",x"60", -- 0x2190
    x"FE",x"8D",x"60",x"FE",x"8E",x"60",x"FE",x"8D", -- 0x2198
    x"60",x"FE",x"8E",x"60",x"FE",x"8D",x"60",x"FE", -- 0x21A0
    x"8E",x"60",x"FE",x"8D",x"60",x"FE",x"8E",x"60", -- 0x21A8
    x"FE",x"8D",x"60",x"FE",x"AD",x"6A",x"FE",x"60", -- 0x21B0
    x"0A",x"2A",x"8D",x"60",x"FE",x"09",x"02",x"8D", -- 0x21B8
    x"60",x"FE",x"2A",x"29",x"FD",x"8D",x"60",x"FE", -- 0x21C0
    x"09",x"02",x"8D",x"60",x"FE",x"2A",x"29",x"FD", -- 0x21C8
    x"8D",x"60",x"FE",x"09",x"02",x"8D",x"60",x"FE", -- 0x21D0
    x"2A",x"29",x"FD",x"8D",x"60",x"FE",x"09",x"02", -- 0x21D8
    x"8D",x"60",x"FE",x"2A",x"29",x"FD",x"8D",x"60", -- 0x21E0
    x"FE",x"09",x"02",x"8D",x"60",x"FE",x"2A",x"29", -- 0x21E8
    x"FD",x"8D",x"60",x"FE",x"09",x"02",x"8D",x"60", -- 0x21F0
    x"FE",x"2A",x"29",x"FD",x"8D",x"60",x"FE",x"09", -- 0x21F8
    x"02",x"8D",x"60",x"FE",x"2A",x"29",x"FD",x"8D", -- 0x2200
    x"60",x"FE",x"09",x"02",x"8D",x"60",x"FE",x"60", -- 0x2208
    x"2C",x"40",x"0D",x"30",x"38",x"A2",x"01",x"A9", -- 0x2210
    x"03",x"8E",x"60",x"FE",x"8D",x"60",x"FE",x"8E", -- 0x2218
    x"60",x"FE",x"8D",x"60",x"FE",x"8E",x"60",x"FE", -- 0x2220
    x"8D",x"60",x"FE",x"8E",x"60",x"FE",x"8D",x"60", -- 0x2228
    x"FE",x"8E",x"60",x"FE",x"8D",x"60",x"FE",x"8E", -- 0x2230
    x"60",x"FE",x"8D",x"60",x"FE",x"8E",x"60",x"FE", -- 0x2238
    x"8D",x"60",x"FE",x"8E",x"60",x"FE",x"8D",x"60", -- 0x2240
    x"FE",x"88",x"D0",x"CD",x"60",x"A9",x"FF",x"8D", -- 0x2248
    x"18",x"FE",x"EA",x"EA",x"EA",x"88",x"D0",x"F7", -- 0x2250
    x"60",x"2C",x"40",x"0D",x"30",x"36",x"8E",x"41", -- 0x2258
    x"0D",x"A0",x"07",x"BD",x"42",x"0D",x"20",x"B8", -- 0x2260
    x"A1",x"E8",x"88",x"D0",x"F6",x"20",x"73",x"A2", -- 0x2268
    x"4C",x"8A",x"A1",x"A9",x"01",x"A2",x"03",x"A0", -- 0x2270
    x"00",x"88",x"F0",x"12",x"8D",x"60",x"FE",x"8E", -- 0x2278
    x"60",x"FE",x"AD",x"6A",x"FE",x"29",x"01",x"D0", -- 0x2280
    x"F0",x"A2",x"01",x"A9",x"03",x"60",x"AD",x"6A", -- 0x2288
    x"FE",x"C9",x"00",x"60",x"8E",x"41",x"0D",x"A0", -- 0x2290
    x"08",x"BD",x"42",x"0D",x"8D",x"18",x"FE",x"EA", -- 0x2298
    x"EA",x"E8",x"88",x"D0",x"F4",x"8D",x"18",x"FE", -- 0x22A0
    x"20",x"58",x"A2",x"AD",x"18",x"FE",x"10",x"E3", -- 0x22A8
    x"88",x"D0",x"F5",x"4C",x"91",x"A2",x"2C",x"40", -- 0x22B0
    x"0D",x"30",x"0A",x"A2",x"01",x"20",x"82",x"A1", -- 0x22B8
    x"C9",x"FE",x"D0",x"F9",x"60",x"A2",x"FF",x"8E", -- 0x22C0
    x"18",x"FE",x"20",x"58",x"A2",x"AD",x"18",x"FE", -- 0x22C8
    x"C9",x"FE",x"D0",x"F3",x"60",x"2C",x"40",x"0D", -- 0x22D0
    x"30",x"15",x"A2",x"01",x"AC",x"D6",x"10",x"D0", -- 0x22D8
    x"09",x"20",x"82",x"A1",x"91",x"A0",x"C8",x"D0", -- 0x22E0
    x"F8",x"60",x"A0",x"00",x"4C",x"2D",x"A3",x"A2", -- 0x22E8
    x"FF",x"8E",x"18",x"FE",x"AC",x"D6",x"10",x"D0", -- 0x22F0
    x"16",x"EA",x"EA",x"EA",x"AD",x"18",x"FE",x"8E", -- 0x22F8
    x"18",x"FE",x"91",x"A0",x"C8",x"C0",x"FF",x"D0", -- 0x2300
    x"F3",x"AD",x"18",x"FE",x"91",x"A0",x"60",x"A0", -- 0x2308
    x"00",x"4C",x"5A",x"A3",x"2C",x"40",x"0D",x"30", -- 0x2310
    x"1E",x"A2",x"01",x"AC",x"D6",x"10",x"D0",x"0B", -- 0x2318
    x"20",x"82",x"A1",x"91",x"A0",x"C8",x"C6",x"A7", -- 0x2320
    x"D0",x"F6",x"60",x"A4",x"A7",x"20",x"82",x"A1", -- 0x2328
    x"8D",x"E5",x"FE",x"88",x"D0",x"F7",x"60",x"A2", -- 0x2330
    x"FF",x"8E",x"18",x"FE",x"AC",x"D6",x"10",x"D0", -- 0x2338
    x"17",x"C6",x"A7",x"F0",x"0D",x"AD",x"18",x"FE", -- 0x2340
    x"8E",x"18",x"FE",x"91",x"A0",x"C8",x"C6",x"A7", -- 0x2348
    x"D0",x"F3",x"AD",x"18",x"FE",x"91",x"A0",x"60", -- 0x2350
    x"A4",x"A7",x"88",x"F0",x"1A",x"EA",x"AD",x"18", -- 0x2358
    x"FE",x"8E",x"18",x"FE",x"8D",x"E5",x"FE",x"20", -- 0x2360
    x"58",x"A2",x"20",x"58",x"A2",x"EA",x"EA",x"EA", -- 0x2368
    x"88",x"D0",x"EA",x"EA",x"EA",x"EA",x"EA",x"AD", -- 0x2370
    x"18",x"FE",x"8D",x"E5",x"FE",x"60",x"2C",x"40", -- 0x2378
    x"0D",x"30",x"0E",x"A0",x"00",x"A2",x"01",x"20", -- 0x2380
    x"82",x"A1",x"99",x"00",x"0E",x"C8",x"D0",x"F7", -- 0x2388
    x"60",x"A0",x"00",x"A2",x"FF",x"8E",x"18",x"FE", -- 0x2390
    x"20",x"58",x"A2",x"AD",x"18",x"FE",x"8E",x"18", -- 0x2398
    x"FE",x"99",x"00",x"0E",x"C8",x"C0",x"FF",x"D0", -- 0x23A0
    x"F2",x"AD",x"18",x"FE",x"99",x"00",x"0E",x"60", -- 0x23A8
    x"2C",x"40",x"0D",x"30",x"0A",x"A0",x"02",x"20", -- 0x23B0
    x"15",x"A2",x"A9",x"FE",x"4C",x"B8",x"A1",x"A2", -- 0x23B8
    x"FF",x"8E",x"18",x"FE",x"20",x"58",x"A2",x"8E", -- 0x23C0
    x"18",x"FE",x"20",x"58",x"A2",x"CA",x"8E",x"18", -- 0x23C8
    x"FE",x"60",x"A0",x"02",x"2C",x"40",x"0D",x"30", -- 0x23D0
    x"1A",x"20",x"15",x"A2",x"20",x"73",x"A2",x"20", -- 0x23D8
    x"9C",x"A1",x"A8",x"29",x"1F",x"C9",x"05",x"D0", -- 0x23E0
    x"2D",x"A2",x"01",x"20",x"82",x"A1",x"C9",x"FF", -- 0x23E8
    x"D0",x"F9",x"60",x"20",x"4D",x"A2",x"A2",x"FF", -- 0x23F0
    x"8E",x"18",x"FE",x"20",x"58",x"A2",x"AD",x"18", -- 0x23F8
    x"FE",x"A8",x"29",x"1F",x"C9",x"05",x"D0",x"0E", -- 0x2400
    x"A9",x"FF",x"8E",x"18",x"FE",x"20",x"58",x"A2", -- 0x2408
    x"CD",x"18",x"FE",x"D0",x"F5",x"60",x"98",x"20", -- 0x2410
    x"1F",x"A0",x"C5",x"4D",x"4D",x"43",x"20",x"57", -- 0x2418
    x"72",x"69",x"74",x"65",x"20",x"72",x"65",x"73", -- 0x2420
    x"70",x"6F",x"6E",x"73",x"65",x"20",x"66",x"61", -- 0x2428
    x"75",x"6C",x"74",x"20",x"00",x"2C",x"40",x"0D", -- 0x2430
    x"30",x"1A",x"AC",x"D6",x"10",x"D0",x"09",x"B1", -- 0x2438
    x"A0",x"20",x"B8",x"A1",x"C8",x"D0",x"F8",x"60", -- 0x2440
    x"A0",x"00",x"AD",x"E5",x"FE",x"20",x"B8",x"A1", -- 0x2448
    x"C8",x"D0",x"F7",x"60",x"AC",x"D6",x"10",x"D0", -- 0x2450
    x"09",x"B1",x"A0",x"8D",x"18",x"FE",x"C8",x"D0", -- 0x2458
    x"F8",x"60",x"A0",x"00",x"AD",x"E5",x"FE",x"8D", -- 0x2460
    x"18",x"FE",x"20",x"58",x"A2",x"20",x"58",x"A2", -- 0x2468
    x"20",x"58",x"A2",x"C8",x"D0",x"EE",x"60",x"2C", -- 0x2470
    x"40",x"0D",x"30",x"0C",x"A0",x"00",x"B9",x"00", -- 0x2478
    x"0E",x"20",x"B8",x"A1",x"C8",x"D0",x"F7",x"60", -- 0x2480
    x"A0",x"00",x"EA",x"B9",x"00",x"0E",x"8D",x"18", -- 0x2488
    x"FE",x"C8",x"D0",x"F6",x"60",x"9D",x"43",x"0D", -- 0x2490
    x"A9",x"00",x"9D",x"44",x"0D",x"9D",x"45",x"0D", -- 0x2498
    x"9D",x"46",x"0D",x"9D",x"47",x"0D",x"A9",x"FF", -- 0x24A0
    x"9D",x"42",x"0D",x"9D",x"48",x"0D",x"9D",x"49", -- 0x24A8
    x"0D",x"AE",x"03",x"0D",x"BD",x"D2",x"A4",x"8D", -- 0x24B0
    x"40",x"0D",x"60",x"2C",x"C9",x"10",x"30",x"11", -- 0x24B8
    x"A9",x"8F",x"A2",x"0C",x"A0",x"FF",x"20",x"F4", -- 0x24C0
    x"FF",x"8C",x"01",x"0D",x"A9",x"FF",x"8D",x"C9", -- 0x24C8
    x"10",x"60",x"80",x"00",x"A9",x"03",x"8D",x"62", -- 0x24D0
    x"FE",x"A9",x"00",x"8D",x"60",x"FE",x"AD",x"6B", -- 0x24D8
    x"FE",x"29",x"E3",x"8D",x"6B",x"FE",x"A9",x"1C", -- 0x24E0
    x"8D",x"6E",x"FE",x"60",x"AD",x"02",x"0D",x"C9", -- 0x24E8
    x"54",x"D0",x"04",x"20",x"D4",x"A4",x"60",x"20", -- 0x24F0
    x"06",x"A5",x"D0",x"FA",x"20",x"00",x"A0",x"FF", -- 0x24F8
    x"43",x"61",x"72",x"64",x"3F",x"00",x"20",x"71", -- 0x2500
    x"A1",x"A2",x"FF",x"8E",x"03",x"0D",x"20",x"BB", -- 0x2508
    x"A4",x"A2",x"00",x"A9",x"40",x"20",x"95",x"A4", -- 0x2510
    x"A9",x"95",x"8D",x"48",x"0D",x"A2",x"08",x"A9", -- 0x2518
    x"41",x"20",x"95",x"A4",x"20",x"D4",x"A4",x"A9", -- 0x2520
    x"32",x"85",x"A6",x"AE",x"04",x"0D",x"E0",x"02", -- 0x2528
    x"B0",x"5A",x"8E",x"03",x"0D",x"BD",x"D2",x"A4", -- 0x2530
    x"8D",x"40",x"0D",x"A0",x"0A",x"20",x"10",x"A2", -- 0x2538
    x"A2",x"00",x"20",x"59",x"A2",x"29",x"81",x"C9", -- 0x2540
    x"01",x"D0",x"35",x"24",x"FF",x"30",x"31",x"A2", -- 0x2548
    x"08",x"20",x"59",x"A2",x"C9",x"02",x"B0",x"28", -- 0x2550
    x"C9",x"00",x"D0",x"EF",x"A2",x"00",x"A9",x"50", -- 0x2558
    x"20",x"95",x"A4",x"A9",x"02",x"8D",x"46",x"0D", -- 0x2560
    x"A2",x"00",x"20",x"59",x"A2",x"D0",x"23",x"A9", -- 0x2568
    x"54",x"8D",x"02",x"0D",x"AD",x"03",x"0D",x"8D", -- 0x2570
    x"04",x"0D",x"20",x"7B",x"A1",x"A9",x"FF",x"60", -- 0x2578
    x"AE",x"03",x"0D",x"E8",x"E0",x"02",x"90",x"AA", -- 0x2580
    x"C6",x"A6",x"D0",x"9F",x"A9",x"00",x"8D",x"02", -- 0x2588
    x"0D",x"60",x"20",x"1F",x"A0",x"FF",x"53",x"65", -- 0x2590
    x"74",x"20",x"62",x"6C",x"6F",x"63",x"6B",x"20", -- 0x2598
    x"6C",x"65",x"6E",x"20",x"65",x"72",x"72",x"6F", -- 0x25A0
    x"72",x"20",x"00",x"A9",x"51",x"A2",x"00",x"20", -- 0x25A8
    x"95",x"A4",x"A5",x"A2",x"8D",x"46",x"0D",x"A5", -- 0x25B0
    x"A3",x"8D",x"45",x"0D",x"A5",x"A4",x"8D",x"44", -- 0x25B8
    x"0D",x"60",x"A2",x"00",x"20",x"59",x"A2",x"D0", -- 0x25C0
    x"04",x"20",x"B6",x"A2",x"60",x"20",x"1F",x"A0", -- 0x25C8
    x"C5",x"4D",x"4D",x"43",x"20",x"52",x"65",x"61", -- 0x25D0
    x"64",x"20",x"66",x"61",x"75",x"6C",x"74",x"20", -- 0x25D8
    x"00",x"A2",x"00",x"20",x"59",x"A2",x"D0",x"03", -- 0x25E0
    x"4C",x"B0",x"A3",x"20",x"1F",x"A0",x"C5",x"4D", -- 0x25E8
    x"4D",x"43",x"20",x"57",x"72",x"69",x"74",x"65", -- 0x25F0
    x"20",x"66",x"61",x"75",x"6C",x"74",x"20",x"00", -- 0x25F8
    x"20",x"71",x"A1",x"A9",x"00",x"8D",x"D6",x"10", -- 0x2600
    x"85",x"A0",x"A9",x"0E",x"85",x"A1",x"60",x"20", -- 0x2608
    x"00",x"A6",x"20",x"AB",x"A5",x"20",x"C2",x"A5", -- 0x2610
    x"20",x"D5",x"A2",x"E6",x"A1",x"20",x"D5",x"A2", -- 0x2618
    x"A0",x"02",x"20",x"10",x"A2",x"4C",x"7B",x"A1", -- 0x2620
    x"20",x"00",x"A6",x"A9",x"58",x"20",x"AD",x"A5", -- 0x2628
    x"20",x"E1",x"A5",x"20",x"35",x"A4",x"E6",x"A1", -- 0x2630
    x"20",x"35",x"A4",x"20",x"D2",x"A3",x"4C",x"7B", -- 0x2638
    x"A1",x"60",x"20",x"71",x"A1",x"20",x"4B",x"A6", -- 0x2640
    x"4C",x"7B",x"A1",x"A6",x"A5",x"F0",x"F2",x"A9", -- 0x2648
    x"01",x"20",x"98",x"A0",x"A6",x"A5",x"66",x"A2", -- 0x2650
    x"66",x"A6",x"10",x"01",x"E8",x"86",x"A5",x"06", -- 0x2658
    x"A2",x"20",x"AB",x"A5",x"A6",x"A5",x"E0",x"03", -- 0x2660
    x"B0",x"08",x"A5",x"A7",x"D0",x"4F",x"E0",x"01", -- 0x2668
    x"F0",x"42",x"24",x"A6",x"10",x"0D",x"20",x"C2", -- 0x2670
    x"A5",x"A0",x"00",x"84",x"A6",x"20",x"10",x"A2", -- 0x2678
    x"4C",x"8B",x"A6",x"20",x"C2",x"A5",x"20",x"D5", -- 0x2680
    x"A2",x"E6",x"A1",x"20",x"D5",x"A2",x"E6",x"A1", -- 0x2688
    x"A0",x"02",x"20",x"10",x"A2",x"EE",x"46",x"0D", -- 0x2690
    x"EE",x"46",x"0D",x"D0",x"08",x"EE",x"45",x"0D", -- 0x2698
    x"D0",x"03",x"EE",x"44",x"0D",x"A6",x"A5",x"CA", -- 0x26A0
    x"CA",x"F0",x"96",x"86",x"A5",x"E0",x"03",x"B0", -- 0x26A8
    x"D2",x"4C",x"6A",x"A6",x"20",x"C2",x"A5",x"20", -- 0x26B0
    x"D5",x"A2",x"4C",x"E4",x"A6",x"20",x"C2",x"A5", -- 0x26B8
    x"24",x"A6",x"10",x"08",x"A0",x"00",x"20",x"10", -- 0x26C0
    x"A2",x"4C",x"D5",x"A6",x"C6",x"A5",x"F0",x"05", -- 0x26C8
    x"20",x"D5",x"A2",x"E6",x"A1",x"20",x"14",x"A3", -- 0x26D0
    x"98",x"49",x"FF",x"A8",x"C8",x"20",x"10",x"A2", -- 0x26D8
    x"A5",x"A5",x"D0",x"05",x"A0",x"00",x"20",x"10", -- 0x26E0
    x"A2",x"A0",x"02",x"4C",x"10",x"A2",x"60",x"20", -- 0x26E8
    x"71",x"A1",x"20",x"F8",x"A6",x"4C",x"7B",x"A1", -- 0x26F0
    x"A6",x"A5",x"F0",x"F2",x"A9",x"00",x"20",x"98", -- 0x26F8
    x"A0",x"A6",x"A5",x"66",x"A2",x"6A",x"06",x"A2", -- 0x2700
    x"48",x"A9",x"58",x"20",x"AD",x"A5",x"68",x"10", -- 0x2708
    x"41",x"A9",x"FF",x"8D",x"82",x"10",x"A9",x"51", -- 0x2710
    x"8D",x"43",x"0D",x"20",x"C2",x"A5",x"20",x"7E", -- 0x2718
    x"A3",x"A0",x"00",x"20",x"10",x"A2",x"A0",x"02", -- 0x2720
    x"20",x"10",x"A2",x"A9",x"58",x"8D",x"43",x"0D", -- 0x2728
    x"20",x"E1",x"A5",x"20",x"77",x"A4",x"20",x"35", -- 0x2730
    x"A4",x"20",x"D2",x"A3",x"C6",x"A5",x"F0",x"AE", -- 0x2738
    x"E6",x"A1",x"EE",x"46",x"0D",x"EE",x"46",x"0D", -- 0x2740
    x"D0",x"08",x"EE",x"45",x"0D",x"D0",x"03",x"EE", -- 0x2748
    x"44",x"0D",x"A6",x"A5",x"F0",x"44",x"CA",x"D0", -- 0x2750
    x"2B",x"A9",x"FF",x"8D",x"82",x"10",x"A9",x"51", -- 0x2758
    x"8D",x"43",x"0D",x"20",x"C2",x"A5",x"A0",x"00", -- 0x2760
    x"20",x"10",x"A2",x"20",x"7E",x"A3",x"A0",x"02", -- 0x2768
    x"20",x"10",x"A2",x"A9",x"58",x"8D",x"43",x"0D", -- 0x2770
    x"20",x"E1",x"A5",x"20",x"35",x"A4",x"20",x"77", -- 0x2778
    x"A4",x"4C",x"D2",x"A3",x"20",x"E1",x"A5",x"20", -- 0x2780
    x"35",x"A4",x"E6",x"A1",x"20",x"35",x"A4",x"E6", -- 0x2788
    x"A1",x"20",x"D2",x"A3",x"C6",x"A5",x"C6",x"A5", -- 0x2790
    x"D0",x"A8",x"60",x"A9",x"51",x"A2",x"08",x"20", -- 0x2798
    x"95",x"A4",x"A5",x"A2",x"8D",x"4E",x"0D",x"A5", -- 0x27A0
    x"A3",x"8D",x"4D",x"0D",x"A5",x"A4",x"8D",x"4C", -- 0x27A8
    x"0D",x"60",x"20",x"71",x"A1",x"A2",x"08",x"20", -- 0x27B0
    x"C4",x"A5",x"A9",x"5F",x"85",x"A0",x"A9",x"0D", -- 0x27B8
    x"85",x"A1",x"A9",x"08",x"85",x"A7",x"20",x"14", -- 0x27C0
    x"A3",x"A0",x"F8",x"20",x"10",x"A2",x"A9",x"67", -- 0x27C8
    x"85",x"A0",x"A9",x"08",x"85",x"A7",x"20",x"14", -- 0x27D0
    x"A3",x"A0",x"FA",x"20",x"10",x"A2",x"18",x"AD", -- 0x27D8
    x"4E",x"0D",x"69",x"20",x"8D",x"4E",x"0D",x"AD", -- 0x27E0
    x"4D",x"0D",x"69",x"03",x"8D",x"4D",x"0D",x"90", -- 0x27E8
    x"03",x"EE",x"4C",x"0D",x"4C",x"7B",x"A1",x"20", -- 0x27F0
    x"06",x"A5",x"F0",x"B5",x"A9",x"7A",x"20",x"F4", -- 0x27F8
    x"FF",x"8A",x"30",x"0D",x"C9",x"65",x"F0",x"04", -- 0x2800
    x"C9",x"42",x"D0",x"A5",x"A9",x"78",x"20",x"F4", -- 0x2808
    x"FF",x"8E",x"52",x"0D",x"4C",x"20",x"93",x"AD", -- 0x2810
    x"05",x"0D",x"C9",x"54",x"D0",x"17",x"AD",x"06", -- 0x2818
    x"0D",x"4D",x"09",x"0D",x"4D",x"07",x"0D",x"4D", -- 0x2820
    x"0A",x"0D",x"4D",x"08",x"0D",x"4D",x"0B",x"0D", -- 0x2828
    x"C9",x"FF",x"D0",x"01",x"60",x"A2",x"08",x"B5", -- 0x2830
    x"A1",x"48",x"CA",x"D0",x"FA",x"A9",x"00",x"85", -- 0x2838
    x"A2",x"85",x"A3",x"85",x"A4",x"20",x"0F",x"A6", -- 0x2840
    x"A9",x"DD",x"8D",x"82",x"10",x"20",x"6B",x"A8", -- 0x2848
    x"F0",x"29",x"A9",x"00",x"8D",x"06",x"0D",x"8D", -- 0x2850
    x"07",x"0D",x"8D",x"08",x"0D",x"A9",x"FF",x"8D", -- 0x2858
    x"09",x"0D",x"8D",x"0A",x"0D",x"8D",x"0B",x"0D", -- 0x2860
    x"4C",x"99",x"A9",x"AD",x"FE",x"0F",x"C9",x"55", -- 0x2868
    x"D0",x"05",x"AD",x"FF",x"0F",x"C9",x"AA",x"60", -- 0x2870
    x"4C",x"A9",x"A9",x"AD",x"C6",x"0F",x"0A",x"85", -- 0x2878
    x"A2",x"AD",x"C7",x"0F",x"2A",x"85",x"A3",x"AD", -- 0x2880
    x"C8",x"0F",x"2A",x"B0",x"EB",x"85",x"A4",x"AD", -- 0x2888
    x"C9",x"0F",x"D0",x"E4",x"20",x"0F",x"A6",x"20", -- 0x2890
    x"6B",x"A8",x"D0",x"DC",x"AD",x"0B",x"0E",x"D0", -- 0x2898
    x"D7",x"AD",x"0C",x"0E",x"C9",x"02",x"D0",x"D0", -- 0x28A0
    x"AD",x"11",x"0E",x"85",x"A5",x"AD",x"12",x"0E", -- 0x28A8
    x"4A",x"66",x"A5",x"4A",x"66",x"A5",x"4A",x"66", -- 0x28B0
    x"A5",x"85",x"A6",x"AD",x"0D",x"0E",x"85",x"A7", -- 0x28B8
    x"AD",x"0E",x"0E",x"0A",x"2E",x"0F",x"0E",x"B0", -- 0x28C0
    x"AF",x"65",x"A2",x"85",x"A2",x"AD",x"0F",x"0E", -- 0x28C8
    x"65",x"A3",x"85",x"A3",x"90",x"02",x"E6",x"A4", -- 0x28D0
    x"0E",x"16",x"0E",x"2E",x"17",x"0E",x"B0",x"98", -- 0x28D8
    x"AE",x"10",x"0E",x"18",x"A5",x"A2",x"6D",x"16", -- 0x28E0
    x"0E",x"85",x"A2",x"A5",x"A3",x"6D",x"17",x"0E", -- 0x28E8
    x"85",x"A3",x"90",x"02",x"E6",x"A4",x"CA",x"D0", -- 0x28F0
    x"EA",x"20",x"0F",x"A6",x"A9",x"00",x"85",x"A8", -- 0x28F8
    x"A9",x"0E",x"85",x"A9",x"A0",x"0B",x"B1",x"A8", -- 0x2900
    x"29",x"0F",x"D0",x"10",x"A0",x"00",x"B1",x"A8", -- 0x2908
    x"D9",x"C2",x"A9",x"D0",x"07",x"C8",x"C0",x"0B", -- 0x2910
    x"F0",x"20",x"D0",x"F2",x"18",x"A5",x"A8",x"69", -- 0x2918
    x"20",x"85",x"A8",x"D0",x"DF",x"20",x"00",x"A0", -- 0x2920
    x"FF",x"49",x"6D",x"61",x"67",x"65",x"20",x"6E", -- 0x2928
    x"6F",x"74",x"20",x"66",x"6F",x"75",x"6E",x"64", -- 0x2930
    x"21",x"00",x"18",x"A5",x"A2",x"65",x"A5",x"85", -- 0x2938
    x"A2",x"A5",x"A3",x"65",x"A6",x"85",x"A3",x"90", -- 0x2940
    x"02",x"E6",x"A4",x"A0",x"1B",x"B1",x"A8",x"48", -- 0x2948
    x"88",x"B1",x"A8",x"38",x"E9",x"02",x"85",x"A8", -- 0x2950
    x"68",x"E9",x"00",x"85",x"A9",x"05",x"A8",x"F0", -- 0x2958
    x"1A",x"06",x"A8",x"26",x"A9",x"A6",x"A7",x"18", -- 0x2960
    x"A5",x"A2",x"65",x"A8",x"85",x"A2",x"A5",x"A3", -- 0x2968
    x"65",x"A9",x"85",x"A3",x"90",x"02",x"E6",x"A4", -- 0x2970
    x"CA",x"D0",x"EC",x"A5",x"A2",x"8D",x"06",x"0D", -- 0x2978
    x"49",x"FF",x"8D",x"09",x"0D",x"A5",x"A3",x"8D", -- 0x2980
    x"07",x"0D",x"49",x"FF",x"8D",x"0A",x"0D",x"A5", -- 0x2988
    x"A4",x"8D",x"08",x"0D",x"49",x"FF",x"8D",x"0B", -- 0x2990
    x"0D",x"A9",x"54",x"8D",x"05",x"0D",x"A2",x"00", -- 0x2998
    x"68",x"95",x"A2",x"E8",x"E0",x"08",x"D0",x"F8", -- 0x29A0
    x"60",x"20",x"00",x"A0",x"FF",x"55",x"6E",x"72", -- 0x29A8
    x"65",x"63",x"6F",x"67",x"6E",x"69",x"73",x"65", -- 0x29B0
    x"64",x"20",x"66",x"6F",x"72",x"6D",x"61",x"74", -- 0x29B8
    x"21",x"00",x"42",x"45",x"45",x"42",x"20",x"20", -- 0x29C0
    x"20",x"20",x"4D",x"4D",x"42",x"08",x"AA",x"20", -- 0x29C8
    x"02",x"AA",x"85",x"B2",x"48",x"20",x"1E",x"AA", -- 0x29D0
    x"8A",x"E5",x"B0",x"AA",x"68",x"20",x"02",x"AA", -- 0x29D8
    x"48",x"20",x"1E",x"AA",x"A5",x"B2",x"E5",x"B0", -- 0x29E0
    x"0A",x"0A",x"0A",x"0A",x"85",x"B2",x"8A",x"05", -- 0x29E8
    x"B2",x"AA",x"68",x"28",x"90",x"0B",x"48",x"8A", -- 0x29F0
    x"F8",x"18",x"69",x"56",x"AA",x"68",x"69",x"02", -- 0x29F8
    x"D8",x"60",x"A0",x"00",x"84",x"B1",x"A0",x"A0", -- 0x2A00
    x"84",x"B0",x"A0",x"05",x"C5",x"B0",x"90",x"04", -- 0x2A08
    x"38",x"E5",x"B0",x"38",x"26",x"B1",x"46",x"B0", -- 0x2A10
    x"88",x"D0",x"F1",x"A5",x"B1",x"60",x"48",x"0A", -- 0x2A18
    x"0A",x"0A",x"85",x"B0",x"68",x"0A",x"18",x"65", -- 0x2A20
    x"B0",x"85",x"B0",x"38",x"60",x"E0",x"FF",x"F0", -- 0x2A28
    x"35",x"BD",x"10",x"0D",x"30",x"30",x"49",x"FF", -- 0x2A30
    x"DD",x"18",x"0D",x"D0",x"24",x"BD",x"0C",x"0D", -- 0x2A38
    x"49",x"FF",x"DD",x"14",x"0D",x"D0",x"1A",x"BD", -- 0x2A40
    x"1C",x"0D",x"C9",x"54",x"F0",x"29",x"20",x"00", -- 0x2A48
    x"A0",x"C9",x"44",x"69",x"73",x"6B",x"20",x"72", -- 0x2A50
    x"65",x"61",x"64",x"20",x"6F",x"6E",x"6C",x"79", -- 0x2A58
    x"00",x"A9",x"FF",x"9D",x"10",x"0D",x"20",x"00", -- 0x2A60
    x"A0",x"C7",x"4E",x"6F",x"20",x"64",x"69",x"73", -- 0x2A68
    x"6B",x"00",x"A9",x"54",x"9D",x"1C",x"0D",x"60", -- 0x2A70
    x"A9",x"00",x"9D",x"1C",x"0D",x"60",x"BD",x"10", -- 0x2A78
    x"0D",x"30",x"E3",x"6A",x"BD",x"0C",x"0D",x"08", -- 0x2A80
    x"AA",x"A9",x"00",x"85",x"A2",x"2A",x"48",x"85", -- 0x2A88
    x"A4",x"8A",x"0A",x"26",x"A4",x"85",x"A3",x"8A", -- 0x2A90
    x"65",x"A3",x"85",x"A3",x"68",x"69",x"00",x"65", -- 0x2A98
    x"A4",x"85",x"A4",x"66",x"A2",x"8A",x"28",x"6A", -- 0x2AA0
    x"66",x"A2",x"4A",x"66",x"A2",x"4A",x"66",x"A2", -- 0x2AA8
    x"65",x"A3",x"85",x"A3",x"A5",x"A4",x"69",x"00", -- 0x2AB0
    x"85",x"A4",x"20",x"17",x"A8",x"38",x"A5",x"A2", -- 0x2AB8
    x"09",x"1F",x"6D",x"06",x"0D",x"85",x"A2",x"A5", -- 0x2AC0
    x"A3",x"6D",x"07",x"0D",x"85",x"A3",x"A5",x"A4", -- 0x2AC8
    x"6D",x"08",x"0D",x"85",x"A4",x"60",x"A5",x"BE", -- 0x2AD0
    x"85",x"A0",x"A5",x"BF",x"85",x"A1",x"A6",x"CF", -- 0x2AD8
    x"20",x"7E",x"AA",x"18",x"A5",x"C5",x"65",x"A2", -- 0x2AE0
    x"85",x"A2",x"A5",x"C4",x"29",x"03",x"48",x"65", -- 0x2AE8
    x"A3",x"85",x"A3",x"90",x"02",x"E6",x"A4",x"A5", -- 0x2AF0
    x"C3",x"85",x"A5",x"A5",x"C4",x"4A",x"4A",x"4A", -- 0x2AF8
    x"4A",x"29",x"03",x"D0",x"1E",x"A5",x"C2",x"85", -- 0x2B00
    x"A7",x"F0",x"04",x"E6",x"A5",x"F0",x"14",x"18", -- 0x2B08
    x"A5",x"C5",x"65",x"A5",x"AA",x"68",x"69",x"00", -- 0x2B10
    x"C9",x"03",x"90",x"06",x"D0",x"17",x"E0",x"21", -- 0x2B18
    x"B0",x"13",x"60",x"20",x"00",x"A0",x"FF",x"42", -- 0x2B20
    x"6C",x"6F",x"63",x"6B",x"20",x"74",x"6F",x"6F", -- 0x2B28
    x"20",x"62",x"69",x"67",x"00",x"20",x"00",x"A0", -- 0x2B30
    x"FF",x"44",x"69",x"73",x"6B",x"20",x"6F",x"76", -- 0x2B38
    x"65",x"72",x"66",x"6C",x"6F",x"77",x"00",x"20", -- 0x2B40
    x"4D",x"83",x"20",x"58",x"83",x"20",x"EC",x"A4", -- 0x2B48
    x"A6",x"CF",x"8E",x"20",x"0D",x"20",x"7E",x"AA", -- 0x2B50
    x"20",x"0F",x"A6",x"A5",x"CF",x"8D",x"82",x"10", -- 0x2B58
    x"60",x"20",x"EC",x"A4",x"A6",x"CF",x"20",x"2D", -- 0x2B60
    x"AA",x"20",x"7E",x"AA",x"4C",x"28",x"A6",x"08", -- 0x2B68
    x"48",x"A0",x"FF",x"8C",x"82",x"10",x"C8",x"98", -- 0x2B70
    x"99",x"00",x"0E",x"99",x"00",x"0F",x"C8",x"D0", -- 0x2B78
    x"F7",x"A9",x"03",x"8D",x"06",x"0F",x"A9",x"20", -- 0x2B80
    x"8D",x"07",x"0F",x"20",x"EC",x"A4",x"68",x"28", -- 0x2B88
    x"20",x"87",x"AA",x"4C",x"28",x"A6",x"20",x"EC", -- 0x2B90
    x"A4",x"20",x"D6",x"AA",x"20",x"42",x"A6",x"20", -- 0x2B98
    x"CD",x"A0",x"A9",x"01",x"60",x"20",x"EC",x"A4", -- 0x2BA0
    x"20",x"D6",x"AA",x"A6",x"CF",x"20",x"2D",x"AA", -- 0x2BA8
    x"20",x"EF",x"A6",x"20",x"CD",x"A0",x"A9",x"01", -- 0x2BB0
    x"60",x"A8",x"C8",x"98",x"D0",x"01",x"38",x"2A", -- 0x2BB8
    x"2A",x"2A",x"2A",x"2A",x"48",x"29",x"1F",x"A8", -- 0x2BC0
    x"68",x"09",x"1F",x"6A",x"60",x"20",x"B9",x"AB", -- 0x2BC8
    x"48",x"8A",x"48",x"98",x"48",x"20",x"98",x"AC", -- 0x2BD0
    x"68",x"6A",x"68",x"AA",x"68",x"A8",x"B0",x"04", -- 0x2BD8
    x"B9",x"00",x"0E",x"60",x"B9",x"00",x"0F",x"60", -- 0x2BE0
    x"08",x"48",x"8D",x"5F",x"0D",x"A9",x"00",x"2A", -- 0x2BE8
    x"8D",x"60",x"0D",x"8E",x"61",x"0D",x"A2",x"03", -- 0x2BF0
    x"EC",x"61",x"0D",x"F0",x"15",x"BD",x"0C",x"0D", -- 0x2BF8
    x"CD",x"5F",x"0D",x"D0",x"0D",x"BD",x"10",x"0D", -- 0x2C00
    x"CD",x"60",x"0D",x"D0",x"05",x"A9",x"FF",x"9D", -- 0x2C08
    x"10",x"0D",x"CA",x"10",x"E3",x"AE",x"61",x"0D", -- 0x2C10
    x"68",x"28",x"60",x"08",x"48",x"9D",x"0C",x"0D", -- 0x2C18
    x"49",x"FF",x"9D",x"14",x"0D",x"A9",x"00",x"2A", -- 0x2C20
    x"9D",x"10",x"0D",x"49",x"FF",x"9D",x"18",x"0D", -- 0x2C28
    x"68",x"28",x"20",x"E8",x"AB",x"20",x"CD",x"AB", -- 0x2C30
    x"30",x"08",x"F0",x"03",x"4C",x"72",x"AA",x"4C", -- 0x2C38
    x"78",x"AA",x"A8",x"A9",x"FF",x"9D",x"10",x"0D", -- 0x2C40
    x"C8",x"D0",x"1A",x"20",x"00",x"A0",x"C7",x"44", -- 0x2C48
    x"69",x"73",x"6B",x"20",x"6E",x"75",x"6D",x"62", -- 0x2C50
    x"65",x"72",x"20",x"6E",x"6F",x"74",x"20",x"76", -- 0x2C58
    x"61",x"6C",x"69",x"64",x"00",x"20",x"00",x"A0", -- 0x2C60
    x"C7",x"44",x"69",x"73",x"6B",x"20",x"6E",x"6F", -- 0x2C68
    x"74",x"20",x"66",x"6F",x"72",x"6D",x"61",x"74", -- 0x2C70
    x"74",x"65",x"64",x"00",x"29",x"7E",x"48",x"20", -- 0x2C78
    x"17",x"A8",x"18",x"68",x"6D",x"06",x"0D",x"85", -- 0x2C80
    x"A2",x"AD",x"07",x"0D",x"69",x"00",x"85",x"A3", -- 0x2C88
    x"AD",x"08",x"0D",x"69",x"00",x"85",x"A4",x"60", -- 0x2C90
    x"29",x"FE",x"09",x"80",x"CD",x"82",x"10",x"F0", -- 0x2C98
    x"F6",x"8D",x"82",x"10",x"48",x"20",x"EC",x"A4", -- 0x2CA0
    x"68",x"20",x"7C",x"AC",x"4C",x"0F",x"A6",x"8D", -- 0x2CA8
    x"82",x"10",x"20",x"7C",x"AC",x"4C",x"0F",x"A6", -- 0x2CB0
    x"20",x"EC",x"A4",x"AD",x"82",x"10",x"20",x"7C", -- 0x2CB8
    x"AC",x"4C",x"28",x"A6",x"AD",x"82",x"10",x"20", -- 0x2CC0
    x"7C",x"AC",x"4C",x"28",x"A6",x"20",x"B8",x"AC", -- 0x2CC8
    x"A2",x"03",x"20",x"D9",x"AC",x"CA",x"10",x"FA", -- 0x2CD0
    x"60",x"BD",x"10",x"0D",x"30",x"2B",x"49",x"FF", -- 0x2CD8
    x"DD",x"18",x"0D",x"D0",x"18",x"BD",x"0C",x"0D", -- 0x2CE0
    x"49",x"FF",x"DD",x"14",x"0D",x"D0",x"0E",x"BD", -- 0x2CE8
    x"10",x"0D",x"6A",x"BD",x"0C",x"0D",x"20",x"CD", -- 0x2CF0
    x"AB",x"F0",x"0B",x"10",x"07",x"A9",x"FF",x"9D", -- 0x2CF8
    x"10",x"0D",x"D0",x"02",x"A9",x"54",x"9D",x"1C", -- 0x2D00
    x"0D",x"60",x"A9",x"FF",x"A2",x"1F",x"9D",x"20", -- 0x2D08
    x"0D",x"CA",x"D0",x"FA",x"8E",x"04",x"0D",x"A9", -- 0x2D10
    x"00",x"8D",x"02",x"0D",x"8D",x"05",x"0D",x"8D", -- 0x2D18
    x"20",x"0D",x"A9",x"80",x"20",x"A1",x"AC",x"A2", -- 0x2D20
    x"00",x"AD",x"52",x"0D",x"C9",x"42",x"F0",x"16", -- 0x2D28
    x"BD",x"10",x"0D",x"30",x"43",x"49",x"FF",x"DD", -- 0x2D30
    x"18",x"0D",x"D0",x"0A",x"BD",x"0C",x"0D",x"49", -- 0x2D38
    x"FF",x"DD",x"14",x"0D",x"F0",x"16",x"BD",x"00", -- 0x2D40
    x"0E",x"9D",x"0C",x"0D",x"49",x"FF",x"9D",x"14", -- 0x2D48
    x"0D",x"BD",x"04",x"0E",x"9D",x"10",x"0D",x"49", -- 0x2D50
    x"FF",x"9D",x"18",x"0D",x"8A",x"F0",x"1E",x"A8", -- 0x2D58
    x"88",x"BD",x"10",x"0D",x"30",x"17",x"D9",x"10", -- 0x2D60
    x"0D",x"D0",x"08",x"BD",x"0C",x"0D",x"D9",x"0C", -- 0x2D68
    x"0D",x"F0",x"05",x"88",x"10",x"EB",x"30",x"05", -- 0x2D70
    x"A9",x"FF",x"9D",x"10",x"0D",x"E8",x"E0",x"04", -- 0x2D78
    x"D0",x"A7",x"4C",x"D0",x"AC",x"08",x"48",x"8D", -- 0x2D80
    x"53",x"0D",x"A9",x"00",x"2A",x"8D",x"54",x"0D", -- 0x2D88
    x"68",x"28",x"08",x"48",x"20",x"CD",x"A9",x"8E", -- 0x2D90
    x"55",x"0D",x"8D",x"56",x"0D",x"68",x"28",x"20", -- 0x2D98
    x"B9",x"AB",x"29",x"F0",x"85",x"F2",x"98",x"29", -- 0x2DA0
    x"01",x"09",x"0E",x"85",x"F3",x"98",x"29",x"FE", -- 0x2DA8
    x"09",x"80",x"8D",x"52",x"0D",x"20",x"9C",x"AC", -- 0x2DB0
    x"4C",x"19",x"AE",x"A9",x"00",x"8D",x"55",x"0D", -- 0x2DB8
    x"8D",x"56",x"0D",x"8D",x"53",x"0D",x"8D",x"54", -- 0x2DC0
    x"0D",x"A9",x"10",x"85",x"F2",x"A9",x"0E",x"85", -- 0x2DC8
    x"F3",x"A9",x"80",x"8D",x"52",x"0D",x"20",x"9C", -- 0x2DD0
    x"AC",x"4C",x"19",x"AE",x"C9",x"FF",x"F0",x"41", -- 0x2DD8
    x"18",x"A5",x"F2",x"69",x"10",x"85",x"F2",x"D0", -- 0x2DE0
    x"18",x"A5",x"F3",x"49",x"01",x"85",x"F3",x"6A", -- 0x2DE8
    x"B0",x"0F",x"AD",x"52",x"0D",x"69",x"02",x"C9", -- 0x2DF0
    x"A0",x"F0",x"26",x"8D",x"52",x"0D",x"20",x"9C", -- 0x2DF8
    x"AC",x"EE",x"53",x"0D",x"D0",x"03",x"EE",x"54", -- 0x2E00
    x"0D",x"F8",x"18",x"AD",x"55",x"0D",x"69",x"01", -- 0x2E08
    x"8D",x"55",x"0D",x"90",x"03",x"EE",x"56",x"0D", -- 0x2E10
    x"D8",x"A0",x"0F",x"B1",x"F2",x"30",x"BD",x"18", -- 0x2E18
    x"60",x"A9",x"FF",x"8D",x"54",x"0D",x"38",x"60", -- 0x2E20
    x"20",x"EC",x"A4",x"A9",x"80",x"8D",x"52",x"0D", -- 0x2E28
    x"20",x"AF",x"AC",x"A9",x"10",x"85",x"F2",x"A9", -- 0x2E30
    x"0E",x"85",x"F3",x"20",x"17",x"A8",x"18",x"AD", -- 0x2E38
    x"06",x"0D",x"69",x"20",x"85",x"A2",x"AD",x"07", -- 0x2E40
    x"0D",x"69",x"00",x"85",x"A3",x"AD",x"08",x"0D", -- 0x2E48
    x"69",x"00",x"85",x"A4",x"20",x"9B",x"A7",x"A0", -- 0x2E50
    x"0F",x"B1",x"F2",x"C9",x"FF",x"F0",x"39",x"20", -- 0x2E58
    x"B2",x"A7",x"A0",x"0B",x"B9",x"5F",x"0D",x"91", -- 0x2E60
    x"F2",x"88",x"10",x"F8",x"18",x"A5",x"F2",x"69", -- 0x2E68
    x"10",x"85",x"F2",x"D0",x"E2",x"A5",x"F3",x"49", -- 0x2E70
    x"01",x"85",x"F3",x"6A",x"B0",x"D9",x"20",x"C4", -- 0x2E78
    x"AC",x"18",x"AD",x"52",x"0D",x"69",x"02",x"C9", -- 0x2E80
    x"A0",x"F0",x"18",x"8D",x"52",x"0D",x"24",x"FF", -- 0x2E88
    x"30",x"12",x"20",x"AF",x"AC",x"4C",x"57",x"AE", -- 0x2E90
    x"A5",x"F2",x"D0",x"04",x"66",x"F3",x"90",x"03", -- 0x2E98
    x"20",x"C4",x"AC",x"60",x"4C",x"82",x"A0",x"A2", -- 0x2EA0
    x"0B",x"A9",x"00",x"20",x"C6",x"88",x"9D",x"5F", -- 0x2EA8
    x"0D",x"CA",x"10",x"F7",x"E8",x"20",x"C5",x"FF", -- 0x2EB0
    x"B0",x"0A",x"20",x"C6",x"88",x"9D",x"5F",x"0D", -- 0x2EB8
    x"E0",x"0B",x"90",x"F0",x"20",x"B4",x"8A",x"AE", -- 0x2EC0
    x"82",x"10",x"BD",x"10",x"0D",x"6A",x"BD",x"0C", -- 0x2EC8
    x"0D",x"20",x"B9",x"AB",x"29",x"F0",x"48",x"98", -- 0x2ED0
    x"48",x"29",x"FE",x"09",x"80",x"20",x"A1",x"AC", -- 0x2ED8
    x"68",x"18",x"29",x"01",x"69",x"0E",x"85",x"F3", -- 0x2EE0
    x"68",x"85",x"F2",x"A0",x"0B",x"B9",x"5F",x"0D", -- 0x2EE8
    x"91",x"F2",x"88",x"10",x"F8",x"4C",x"B8",x"AC", -- 0x2EF0
    x"44",x"49",x"4E",x"B3",x"C0",x"12",x"44",x"42", -- 0x2EF8
    x"4F",x"4F",x"54",x"B3",x"B5",x"02",x"44",x"43", -- 0x2F00
    x"41",x"54",x"B3",x"C6",x"04",x"44",x"44",x"49", -- 0x2F08
    x"53",x"4B",x"53",x"B5",x"76",x"01",x"44",x"4C", -- 0x2F10
    x"4F",x"43",x"4B",x"B5",x"BC",x"02",x"44",x"55", -- 0x2F18
    x"4E",x"4C",x"4F",x"43",x"4B",x"B5",x"C0",x"02", -- 0x2F20
    x"44",x"46",x"52",x"45",x"45",x"B4",x"B0",x"00", -- 0x2F28
    x"44",x"4B",x"49",x"4C",x"4C",x"B5",x"E3",x"03", -- 0x2F30
    x"44",x"52",x"45",x"53",x"54",x"4F",x"52",x"45", -- 0x2F38
    x"B6",x"26",x"03",x"44",x"4E",x"45",x"57",x"B6", -- 0x2F40
    x"7B",x"01",x"44",x"46",x"4F",x"52",x"4D",x"B6", -- 0x2F48
    x"1E",x"03",x"44",x"4F",x"4E",x"42",x"4F",x"4F", -- 0x2F50
    x"54",x"B7",x"49",x"52",x"44",x"52",x"45",x"43", -- 0x2F58
    x"41",x"54",x"AE",x"27",x"00",x"44",x"52",x"4F", -- 0x2F60
    x"4D",x"B7",x"B0",x"86",x"44",x"4D",x"4F",x"44", -- 0x2F68
    x"45",x"B7",x"64",x"07",x"44",x"53",x"57",x"41", -- 0x2F70
    x"50",x"B7",x"9A",x"00",x"44",x"41",x"42",x"4F", -- 0x2F78
    x"55",x"54",x"AF",x"FA",x"00",x"87",x"D6",x"00", -- 0x2F80
    x"44",x"55",x"54",x"49",x"4C",x"53",x"AF",x"CB", -- 0x2F88
    x"00",x"AF",x"BD",x"00",x"A2",x"A0",x"B1",x"F2", -- 0x2F90
    x"C9",x"0D",x"D0",x"16",x"98",x"E8",x"A0",x"02", -- 0x2F98
    x"20",x"CB",x"99",x"20",x"FF",x"B1",x"20",x"20", -- 0x2FA0
    x"44",x"55",x"54",x"49",x"4C",x"53",x"00",x"4C", -- 0x2FA8
    x"E7",x"FF",x"98",x"48",x"20",x"71",x"86",x"68", -- 0x2FB0
    x"A8",x"A2",x"8D",x"4C",x"29",x"B0",x"C8",x"B1", -- 0x2FB8
    x"F2",x"C9",x"0D",x"F0",x"06",x"C9",x"20",x"F0", -- 0x2FC0
    x"F0",x"D0",x"F3",x"60",x"20",x"E7",x"FF",x"20", -- 0x2FC8
    x"FF",x"B1",x"44",x"46",x"53",x"20",x"30",x"2E", -- 0x2FD0
    x"39",x"30",x"00",x"20",x"E7",x"FF",x"A2",x"00", -- 0x2FD8
    x"A9",x"0E",x"86",x"B5",x"85",x"BF",x"A2",x"00", -- 0x2FE0
    x"A9",x"20",x"20",x"EE",x"FF",x"20",x"EE",x"FF", -- 0x2FE8
    x"20",x"C3",x"B2",x"20",x"E7",x"FF",x"C6",x"BF", -- 0x2FF0
    x"D0",x"EE",x"60",x"20",x"FF",x"B1",x"44",x"55", -- 0x2FF8
    x"54",x"49",x"4C",x"53",x"20",x"62",x"79",x"20", -- 0x3000
    x"4D",x"61",x"72",x"74",x"69",x"6E",x"20",x"4D", -- 0x3008
    x"61",x"74",x"68",x"65",x"72",x"20",x"28",x"31", -- 0x3010
    x"39",x"20",x"4E",x"6F",x"76",x"20",x"32",x"30", -- 0x3018
    x"30",x"38",x"29",x"00",x"4C",x"E7",x"FF",x"A2", -- 0x3020
    x"FD",x"98",x"48",x"E8",x"E8",x"68",x"48",x"A8", -- 0x3028
    x"20",x"6B",x"B0",x"E8",x"BD",x"F8",x"AE",x"30", -- 0x3030
    x"28",x"86",x"B5",x"CA",x"88",x"E8",x"C8",x"BD", -- 0x3038
    x"F8",x"AE",x"30",x"16",x"51",x"F2",x"29",x"5F", -- 0x3040
    x"F0",x"F3",x"CA",x"E8",x"BD",x"F8",x"AE",x"10", -- 0x3048
    x"FA",x"B1",x"F2",x"C9",x"2E",x"D0",x"D4",x"C8", -- 0x3050
    x"B0",x"07",x"B1",x"F2",x"20",x"EE",x"82",x"90", -- 0x3058
    x"CA",x"68",x"BD",x"F8",x"AE",x"48",x"BD",x"F9", -- 0x3060
    x"AE",x"48",x"60",x"B1",x"F2",x"C9",x"0D",x"F0", -- 0x3068
    x"08",x"C8",x"F0",x"07",x"C9",x"20",x"F0",x"F3", -- 0x3070
    x"18",x"88",x"60",x"4C",x"B0",x"B2",x"98",x"48", -- 0x3078
    x"A9",x"00",x"8D",x"55",x"0D",x"8D",x"56",x"0D", -- 0x3080
    x"20",x"6B",x"B0",x"B0",x"62",x"B1",x"F2",x"C9", -- 0x3088
    x"0D",x"F0",x"5C",x"38",x"E9",x"30",x"30",x"57", -- 0x3090
    x"C9",x"0A",x"B0",x"53",x"48",x"AD",x"55",x"0D", -- 0x3098
    x"0A",x"48",x"2E",x"56",x"0D",x"AE",x"56",x"0D", -- 0x30A0
    x"0A",x"2E",x"56",x"0D",x"0A",x"2E",x"56",x"0D", -- 0x30A8
    x"8D",x"55",x"0D",x"68",x"6D",x"55",x"0D",x"8D", -- 0x30B0
    x"55",x"0D",x"8A",x"6D",x"56",x"0D",x"AA",x"68", -- 0x30B8
    x"6D",x"55",x"0D",x"8D",x"55",x"0D",x"8A",x"69", -- 0x30C0
    x"00",x"8D",x"56",x"0D",x"C9",x"02",x"B0",x"1F", -- 0x30C8
    x"C8",x"F0",x"1C",x"B1",x"F2",x"C9",x"0D",x"F0", -- 0x30D0
    x"04",x"C9",x"20",x"D0",x"B6",x"AE",x"55",x"0D", -- 0x30D8
    x"AD",x"56",x"0D",x"F0",x"04",x"E8",x"F0",x"07", -- 0x30E0
    x"CA",x"68",x"AD",x"56",x"0D",x"18",x"60",x"68", -- 0x30E8
    x"A8",x"A9",x"00",x"AA",x"38",x"60",x"A9",x"0D", -- 0x30F0
    x"8D",x"5D",x"0D",x"A2",x"00",x"8E",x"5E",x"0D", -- 0x30F8
    x"20",x"6B",x"B0",x"B0",x"49",x"C9",x"22",x"D0", -- 0x3100
    x"04",x"C8",x"8D",x"5D",x"0D",x"B1",x"F2",x"C9", -- 0x3108
    x"0D",x"F0",x"2C",x"C9",x"20",x"D0",x"0B",x"90", -- 0x3110
    x"52",x"AD",x"5D",x"0D",x"C9",x"22",x"D0",x"28", -- 0x3118
    x"A9",x"20",x"C9",x"22",x"F0",x"19",x"C9",x"2A", -- 0x3120
    x"F0",x"31",x"C9",x"61",x"90",x"06",x"C9",x"7B", -- 0x3128
    x"B0",x"02",x"49",x"20",x"9D",x"5F",x"0D",x"C8", -- 0x3130
    x"E8",x"E0",x"0C",x"D0",x"D0",x"B1",x"F2",x"CD", -- 0x3138
    x"5D",x"0D",x"D0",x"27",x"C9",x"0D",x"F0",x"06", -- 0x3140
    x"C8",x"20",x"6B",x"B0",x"90",x"1D",x"8E",x"5C", -- 0x3148
    x"0D",x"E0",x"0C",x"F0",x"05",x"A9",x"00",x"9D", -- 0x3150
    x"5F",x"0D",x"60",x"8D",x"5E",x"0D",x"AD",x"5D", -- 0x3158
    x"0D",x"C9",x"0D",x"F0",x"E3",x"C8",x"B1",x"F2", -- 0x3160
    x"4C",x"3F",x"B1",x"4C",x"B0",x"B2",x"A0",x"00", -- 0x3168
    x"AE",x"5C",x"0D",x"F0",x"17",x"B1",x"F2",x"F0", -- 0x3170
    x"25",x"C9",x"61",x"90",x"06",x"C9",x"7B",x"B0", -- 0x3178
    x"02",x"49",x"20",x"D9",x"5F",x"0D",x"D0",x"16", -- 0x3180
    x"C8",x"CA",x"D0",x"E9",x"B1",x"F2",x"F0",x"0C", -- 0x3188
    x"AD",x"5C",x"0D",x"C9",x"0C",x"F0",x"05",x"AD", -- 0x3190
    x"5E",x"0D",x"F0",x"02",x"18",x"60",x"38",x"60", -- 0x3198
    x"B0",x"05",x"A9",x"20",x"20",x"EE",x"FF",x"A2", -- 0x31A0
    x"20",x"A0",x"04",x"AD",x"56",x"0D",x"20",x"E1", -- 0x31A8
    x"B1",x"AD",x"55",x"0D",x"20",x"E1",x"B1",x"A9", -- 0x31B0
    x"20",x"20",x"EE",x"FF",x"A0",x"00",x"B1",x"F2", -- 0x31B8
    x"F0",x"08",x"20",x"EE",x"FF",x"C8",x"C0",x"0C", -- 0x31C0
    x"D0",x"F4",x"A9",x"20",x"20",x"EE",x"FF",x"C8", -- 0x31C8
    x"C0",x"0D",x"D0",x"F8",x"AA",x"A0",x"0F",x"B1", -- 0x31D0
    x"F2",x"D0",x"02",x"A2",x"50",x"8A",x"4C",x"EE", -- 0x31D8
    x"FF",x"48",x"4A",x"4A",x"4A",x"4A",x"20",x"EA", -- 0x31E0
    x"B1",x"68",x"29",x"0F",x"F0",x"08",x"A2",x"30", -- 0x31E8
    x"18",x"69",x"30",x"4C",x"EE",x"FF",x"88",x"D0", -- 0x31F0
    x"02",x"A2",x"30",x"8A",x"4C",x"EE",x"FF",x"A2", -- 0x31F8
    x"00",x"68",x"85",x"A0",x"68",x"85",x"A1",x"A0", -- 0x3200
    x"00",x"F0",x"07",x"B1",x"A0",x"F0",x"0B",x"20", -- 0x3208
    x"21",x"B2",x"E6",x"A0",x"D0",x"F5",x"E6",x"A1", -- 0x3210
    x"D0",x"F1",x"A5",x"A1",x"48",x"A5",x"A0",x"48", -- 0x3218
    x"60",x"E0",x"00",x"D0",x"03",x"4C",x"EE",x"FF", -- 0x3220
    x"9D",x"00",x"01",x"E8",x"60",x"08",x"10",x"1C", -- 0x3228
    x"22",x"43",x"49",x"4F",x"58",x"28",x"3C",x"64", -- 0x3230
    x"72",x"76",x"3E",x"29",x"00",x"3C",x"64",x"6E", -- 0x3238
    x"6F",x"3E",x"2F",x"3C",x"64",x"73",x"70",x"3E", -- 0x3240
    x"00",x"3C",x"64",x"6E",x"6F",x"3E",x"00",x"28", -- 0x3248
    x"28",x"3C",x"66",x"72",x"6F",x"6D",x"20",x"64", -- 0x3250
    x"6E",x"6F",x"3E",x"29",x"20",x"3C",x"74",x"6F", -- 0x3258
    x"20",x"64",x"6E",x"6F",x"3E",x"29",x"20",x"28", -- 0x3260
    x"3C",x"61",x"64",x"73",x"70",x"3E",x"29",x"00", -- 0x3268
    x"3C",x"64",x"72",x"76",x"3E",x"00",x"3C",x"66", -- 0x3270
    x"73",x"70",x"3E",x"00",x"28",x"3C",x"6D",x"6F", -- 0x3278
    x"64",x"65",x"3E",x"29",x"00",x"28",x"3C",x"72", -- 0x3280
    x"6F",x"6D",x"3E",x"29",x"00",x"48",x"4A",x"4A", -- 0x3288
    x"4A",x"4A",x"20",x"98",x"B2",x"68",x"29",x"0F", -- 0x3290
    x"A8",x"F0",x"14",x"A9",x"20",x"20",x"21",x"B2", -- 0x3298
    x"B9",x"2C",x"B2",x"A8",x"B9",x"2D",x"B2",x"F0", -- 0x32A0
    x"06",x"20",x"21",x"B2",x"C8",x"D0",x"F5",x"60", -- 0x32A8
    x"A2",x"00",x"8E",x"00",x"01",x"E8",x"20",x"01", -- 0x32B0
    x"B2",x"1A",x"53",x"79",x"6E",x"74",x"61",x"78", -- 0x32B8
    x"3A",x"20",x"00",x"A4",x"B5",x"B9",x"F8",x"AE", -- 0x32C0
    x"30",x"06",x"20",x"21",x"B2",x"C8",x"D0",x"F5", -- 0x32C8
    x"C8",x"C8",x"B9",x"F8",x"AE",x"C8",x"84",x"B5", -- 0x32D0
    x"20",x"8D",x"B2",x"E0",x"00",x"F0",x"08",x"A9", -- 0x32D8
    x"00",x"9D",x"00",x"01",x"4C",x"00",x"01",x"60", -- 0x32E0
    x"4C",x"B0",x"B2",x"20",x"6B",x"B0",x"B0",x"17", -- 0x32E8
    x"20",x"7E",x"B0",x"B0",x"BB",x"48",x"20",x"6B", -- 0x32F0
    x"B0",x"68",x"90",x"B4",x"D0",x"26",x"8A",x"8D", -- 0x32F8
    x"5B",x"0D",x"C9",x"04",x"B0",x"1E",x"60",x"A5", -- 0x3300
    x"CF",x"60",x"20",x"6B",x"B0",x"B0",x"A1",x"20", -- 0x3308
    x"7E",x"B0",x"B0",x"9C",x"48",x"20",x"6B",x"B0", -- 0x3310
    x"68",x"90",x"95",x"60",x"20",x"6B",x"B0",x"B0", -- 0x3318
    x"8F",x"4C",x"75",x"B3",x"20",x"00",x"A0",x"CD", -- 0x3320
    x"42",x"61",x"64",x"20",x"64",x"72",x"69",x"76", -- 0x3328
    x"65",x"00",x"20",x"00",x"A0",x"D6",x"44",x"69", -- 0x3330
    x"73",x"6B",x"20",x"6E",x"6F",x"74",x"20",x"66", -- 0x3338
    x"6F",x"75",x"6E",x"64",x"00",x"20",x"6B",x"B0", -- 0x3340
    x"B0",x"9E",x"A9",x"FF",x"20",x"5D",x"B3",x"08", -- 0x3348
    x"E0",x"04",x"B0",x"33",x"28",x"60",x"20",x"6B", -- 0x3350
    x"B0",x"B0",x"8D",x"A5",x"CF",x"8D",x"5B",x"0D", -- 0x3358
    x"20",x"7E",x"B0",x"B0",x"26",x"48",x"20",x"6B", -- 0x3360
    x"B0",x"B0",x"15",x"68",x"D0",x"B6",x"E0",x"04", -- 0x3368
    x"B0",x"B2",x"8E",x"5B",x"0D",x"20",x"7E",x"B0", -- 0x3370
    x"B0",x"11",x"48",x"20",x"6B",x"B0",x"90",x"07", -- 0x3378
    x"68",x"6A",x"8A",x"AE",x"5B",x"0D",x"60",x"68", -- 0x3380
    x"4C",x"B0",x"B2",x"20",x"F6",x"B0",x"20",x"BB", -- 0x3388
    x"AD",x"AD",x"5C",x"0D",x"F0",x"F2",x"AD",x"5E", -- 0x3390
    x"0D",x"D0",x"ED",x"AD",x"54",x"0D",x"30",x"92", -- 0x3398
    x"20",x"6E",x"B1",x"90",x"06",x"20",x"E0",x"AD", -- 0x33A0
    x"4C",x"9B",x"B3",x"AD",x"54",x"0D",x"6A",x"AD", -- 0x33A8
    x"53",x"0D",x"AE",x"5B",x"0D",x"60",x"20",x"1C", -- 0x33B0
    x"B3",x"A6",x"CF",x"20",x"1B",x"AC",x"4C",x"07", -- 0x33B8
    x"94",x"20",x"56",x"B3",x"4C",x"1B",x"AC",x"A9", -- 0x33C0
    x"00",x"8D",x"57",x"0D",x"8D",x"58",x"0D",x"20", -- 0x33C8
    x"7E",x"B0",x"B0",x"2D",x"8E",x"59",x"0D",x"8E", -- 0x33D0
    x"53",x"0D",x"8D",x"5A",x"0D",x"8D",x"54",x"0D", -- 0x33D8
    x"20",x"7E",x"B0",x"B0",x"25",x"8E",x"59",x"0D", -- 0x33E0
    x"8D",x"5A",x"0D",x"EC",x"53",x"0D",x"ED",x"54", -- 0x33E8
    x"0D",x"10",x"1F",x"20",x"00",x"A0",x"FF",x"42", -- 0x33F0
    x"61",x"64",x"20",x"72",x"61",x"6E",x"67",x"65", -- 0x33F8
    x"00",x"A2",x"FE",x"8E",x"59",x"0D",x"E8",x"8E", -- 0x3400
    x"5A",x"0D",x"A9",x"00",x"8D",x"53",x"0D",x"8D", -- 0x3408
    x"54",x"0D",x"EE",x"59",x"0D",x"D0",x"03",x"EE", -- 0x3410
    x"5A",x"0D",x"20",x"F6",x"B0",x"AD",x"54",x"0D", -- 0x3418
    x"6A",x"AD",x"53",x"0D",x"20",x"85",x"AD",x"A2", -- 0x3420
    x"00",x"AD",x"5C",x"0D",x"D0",x"04",x"CA",x"8E", -- 0x3428
    x"5E",x"0D",x"AD",x"54",x"0D",x"30",x"33",x"AD", -- 0x3430
    x"53",x"0D",x"CD",x"59",x"0D",x"AD",x"54",x"0D", -- 0x3438
    x"ED",x"5A",x"0D",x"B0",x"25",x"20",x"6E",x"B1", -- 0x3440
    x"B0",x"16",x"20",x"A0",x"B1",x"F8",x"18",x"AD", -- 0x3448
    x"57",x"0D",x"69",x"01",x"8D",x"57",x"0D",x"AD", -- 0x3450
    x"58",x"0D",x"69",x"00",x"8D",x"58",x"0D",x"D8", -- 0x3458
    x"24",x"FF",x"30",x"47",x"20",x"E0",x"AD",x"4C", -- 0x3460
    x"32",x"B4",x"A9",x"86",x"20",x"F4",x"FF",x"E0", -- 0x3468
    x"00",x"F0",x"03",x"20",x"E7",x"FF",x"AD",x"58", -- 0x3470
    x"0D",x"A2",x"00",x"A0",x"04",x"20",x"E1",x"B1", -- 0x3478
    x"AD",x"57",x"0D",x"20",x"E1",x"B1",x"20",x"FF", -- 0x3480
    x"B1",x"20",x"64",x"69",x"73",x"6B",x"00",x"AD", -- 0x3488
    x"58",x"0D",x"D0",x"05",x"CE",x"57",x"0D",x"F0", -- 0x3490
    x"05",x"A9",x"73",x"20",x"EE",x"FF",x"20",x"FF", -- 0x3498
    x"B1",x"20",x"66",x"6F",x"75",x"6E",x"64",x"00", -- 0x34A0
    x"4C",x"E7",x"FF",x"4C",x"82",x"A0",x"4C",x"B0", -- 0x34A8
    x"B2",x"20",x"6B",x"B0",x"90",x"F8",x"A2",x"00", -- 0x34B0
    x"8E",x"57",x"0D",x"8E",x"58",x"0D",x"8E",x"59", -- 0x34B8
    x"0D",x"8E",x"5A",x"0D",x"A9",x"80",x"20",x"9C", -- 0x34C0
    x"AC",x"A9",x"10",x"85",x"F2",x"A9",x"0E",x"85", -- 0x34C8
    x"F3",x"A0",x"0F",x"B1",x"F2",x"C9",x"FF",x"F0", -- 0x34D0
    x"42",x"F8",x"A8",x"10",x"0E",x"18",x"AD",x"57", -- 0x34D8
    x"0D",x"69",x"01",x"8D",x"57",x"0D",x"90",x"03", -- 0x34E0
    x"EE",x"58",x"0D",x"18",x"AD",x"59",x"0D",x"69", -- 0x34E8
    x"01",x"8D",x"59",x"0D",x"90",x"03",x"EE",x"5A", -- 0x34F0
    x"0D",x"D8",x"18",x"A5",x"F2",x"69",x"10",x"85", -- 0x34F8
    x"F2",x"D0",x"CE",x"A5",x"F3",x"49",x"01",x"85", -- 0x3500
    x"F3",x"6A",x"B0",x"C5",x"AD",x"82",x"10",x"69", -- 0x3508
    x"02",x"C9",x"A0",x"F0",x"06",x"20",x"9C",x"AC", -- 0x3510
    x"4C",x"D1",x"B4",x"A0",x"04",x"A2",x"00",x"AD", -- 0x3518
    x"58",x"0D",x"20",x"E1",x"B1",x"AD",x"57",x"0D", -- 0x3520
    x"20",x"E1",x"B1",x"20",x"FF",x"B1",x"20",x"6F", -- 0x3528
    x"66",x"20",x"00",x"A2",x"00",x"A0",x"04",x"AD", -- 0x3530
    x"5A",x"0D",x"20",x"E1",x"B1",x"AD",x"59",x"0D", -- 0x3538
    x"20",x"E1",x"B1",x"20",x"FF",x"B1",x"20",x"64", -- 0x3540
    x"69",x"73",x"6B",x"00",x"AD",x"5A",x"0D",x"D0", -- 0x3548
    x"07",x"AD",x"59",x"0D",x"C9",x"01",x"F0",x"05", -- 0x3550
    x"A9",x"73",x"20",x"EE",x"FF",x"20",x"FF",x"B1", -- 0x3558
    x"20",x"66",x"72",x"65",x"65",x"20",x"28",x"75", -- 0x3560
    x"6E",x"66",x"6F",x"72",x"6D",x"61",x"74",x"74", -- 0x3568
    x"65",x"64",x"29",x"00",x"4C",x"E7",x"FF",x"20", -- 0x3570
    x"EB",x"B2",x"A2",x"04",x"8E",x"5B",x"0D",x"A2", -- 0x3578
    x"00",x"B0",x"06",x"AA",x"E8",x"8E",x"5B",x"0D", -- 0x3580
    x"CA",x"8A",x"48",x"A2",x"20",x"A0",x"02",x"20", -- 0x3588
    x"E1",x"B1",x"A9",x"3A",x"20",x"EE",x"FF",x"68", -- 0x3590
    x"AA",x"48",x"BD",x"10",x"0D",x"30",x"0F",x"6A", -- 0x3598
    x"BD",x"0C",x"0D",x"20",x"85",x"AD",x"C9",x"FF", -- 0x35A0
    x"F0",x"04",x"38",x"20",x"A0",x"B1",x"20",x"E7", -- 0x35A8
    x"FF",x"68",x"AA",x"E8",x"EC",x"5B",x"0D",x"90", -- 0x35B0
    x"D0",x"60",x"4C",x"B0",x"B2",x"A9",x"00",x"F0", -- 0x35B8
    x"02",x"A9",x"0F",x"48",x"20",x"1C",x"B3",x"20", -- 0x35C0
    x"CD",x"AB",x"30",x"0E",x"68",x"B0",x"05",x"99", -- 0x35C8
    x"00",x"0E",x"90",x"03",x"99",x"00",x"0F",x"4C", -- 0x35D0
    x"CD",x"AC",x"C9",x"FF",x"F0",x"03",x"4C",x"65", -- 0x35D8
    x"AC",x"4C",x"4B",x"AC",x"20",x"BD",x"9B",x"20", -- 0x35E0
    x"0A",x"B3",x"6A",x"08",x"8A",x"48",x"20",x"CD", -- 0x35E8
    x"AB",x"30",x"E7",x"68",x"28",x"20",x"85",x"AD", -- 0x35F0
    x"20",x"FF",x"B1",x"4B",x"69",x"6C",x"6C",x"00", -- 0x35F8
    x"38",x"20",x"A0",x"B1",x"20",x"FF",x"B1",x"20", -- 0x3600
    x"3A",x"20",x"00",x"20",x"9E",x"9C",x"08",x"20", -- 0x3608
    x"E7",x"FF",x"28",x"D0",x"09",x"A0",x"0F",x"A9", -- 0x3610
    x"F0",x"91",x"F2",x"4C",x"CD",x"AC",x"60",x"A9", -- 0x3618
    x"00",x"20",x"29",x"B6",x"4C",x"6F",x"AB",x"A9", -- 0x3620
    x"01",x"8D",x"5F",x"0D",x"20",x"0A",x"B3",x"6A", -- 0x3628
    x"08",x"8A",x"48",x"20",x"CD",x"AB",x"10",x"26", -- 0x3630
    x"AA",x"E8",x"F0",x"3D",x"98",x"29",x"F0",x"85", -- 0x3638
    x"F2",x"A0",x"0E",x"90",x"01",x"C8",x"84",x"F3", -- 0x3640
    x"A0",x"0F",x"98",x"91",x"F2",x"AD",x"5F",x"0D", -- 0x3648
    x"D0",x"06",x"88",x"91",x"F2",x"88",x"10",x"FB", -- 0x3650
    x"20",x"CD",x"AC",x"68",x"28",x"60",x"20",x"00", -- 0x3658
    x"A0",x"FF",x"44",x"69",x"73",x"6B",x"20",x"61", -- 0x3660
    x"6C",x"72",x"65",x"61",x"64",x"79",x"20",x"66", -- 0x3668
    x"6F",x"72",x"6D",x"61",x"74",x"74",x"65",x"64", -- 0x3670
    x"00",x"4C",x"4B",x"AC",x"20",x"EB",x"B2",x"8D", -- 0x3678
    x"5B",x"0D",x"20",x"E0",x"B6",x"08",x"48",x"A9", -- 0x3680
    x"0F",x"91",x"F2",x"88",x"A9",x"00",x"91",x"F2", -- 0x3688
    x"88",x"10",x"FB",x"20",x"B8",x"AC",x"68",x"28", -- 0x3690
    x"08",x"48",x"20",x"6F",x"AB",x"68",x"28",x"08", -- 0x3698
    x"48",x"AE",x"5B",x"0D",x"20",x"1B",x"AC",x"20", -- 0x36A0
    x"FF",x"B1",x"44",x"69",x"73",x"6B",x"20",x"00", -- 0x36A8
    x"68",x"28",x"20",x"CD",x"A9",x"8E",x"55",x"0D", -- 0x36B0
    x"A2",x"00",x"A0",x"04",x"20",x"E1",x"B1",x"AD", -- 0x36B8
    x"55",x"0D",x"20",x"E1",x"B1",x"20",x"FF",x"B1", -- 0x36C0
    x"20",x"69",x"6E",x"20",x"64",x"72",x"69",x"76", -- 0x36C8
    x"65",x"20",x"00",x"AD",x"5B",x"0D",x"A2",x"00", -- 0x36D0
    x"A0",x"02",x"20",x"E1",x"B1",x"4C",x"E7",x"FF", -- 0x36D8
    x"A9",x"10",x"85",x"F2",x"A9",x"0E",x"85",x"F3", -- 0x36E0
    x"A9",x"80",x"8D",x"52",x"0D",x"20",x"A1",x"AC", -- 0x36E8
    x"A9",x"00",x"8D",x"53",x"0D",x"8D",x"54",x"0D", -- 0x36F0
    x"A0",x"0F",x"B1",x"F2",x"10",x"0C",x"C9",x"FF", -- 0x36F8
    x"F0",x"36",x"AD",x"54",x"0D",x"6A",x"AD",x"53", -- 0x3700
    x"0D",x"60",x"EE",x"53",x"0D",x"D0",x"03",x"EE", -- 0x3708
    x"54",x"0D",x"18",x"A5",x"F2",x"69",x"10",x"85", -- 0x3710
    x"F2",x"D0",x"DF",x"A5",x"F3",x"49",x"01",x"85", -- 0x3718
    x"F3",x"29",x"01",x"D0",x"D5",x"18",x"AD",x"52", -- 0x3720
    x"0D",x"69",x"02",x"C9",x"A0",x"F0",x"09",x"8D", -- 0x3728
    x"52",x"0D",x"20",x"A1",x"AC",x"4C",x"F8",x"B6", -- 0x3730
    x"20",x"00",x"A0",x"FF",x"4E",x"6F",x"20",x"66", -- 0x3738
    x"72",x"65",x"65",x"20",x"64",x"69",x"73",x"6B", -- 0x3740
    x"73",x"00",x"20",x"45",x"B3",x"08",x"48",x"8A", -- 0x3748
    x"48",x"A9",x"80",x"20",x"A1",x"AC",x"68",x"AA", -- 0x3750
    x"68",x"9D",x"00",x"0E",x"68",x"29",x"01",x"9D", -- 0x3758
    x"04",x"0E",x"4C",x"B8",x"AC",x"20",x"6B",x"B0", -- 0x3760
    x"A2",x"00",x"B0",x"0B",x"20",x"7E",x"B0",x"B0", -- 0x3768
    x"16",x"C9",x"00",x"F0",x"02",x"A2",x"01",x"8E", -- 0x3770
    x"04",x"0D",x"20",x"E2",x"8D",x"A2",x"FF",x"A9", -- 0x3778
    x"61",x"8D",x"52",x"0D",x"4C",x"17",x"AD",x"20", -- 0x3780
    x"00",x"A0",x"FF",x"42",x"61",x"64",x"20",x"64", -- 0x3788
    x"72",x"69",x"76",x"65",x"72",x"20",x"6D",x"6F", -- 0x3790
    x"64",x"65",x"00",x"A2",x"1E",x"BC",x"02",x"0D", -- 0x3798
    x"BD",x"21",x"0D",x"9D",x"02",x"0D",x"98",x"9D", -- 0x37A0
    x"21",x"0D",x"CA",x"10",x"F0",x"8E",x"82",x"10", -- 0x37A8
    x"60",x"A9",x"00",x"85",x"A6",x"20",x"C2",x"FF", -- 0x37B0
    x"F0",x"6B",x"B1",x"F2",x"C8",x"C9",x"20",x"F0", -- 0x37B8
    x"F9",x"B1",x"F2",x"88",x"C9",x"20",x"D0",x"23", -- 0x37C0
    x"B1",x"F2",x"38",x"E9",x"30",x"30",x"1C",x"C9", -- 0x37C8
    x"0A",x"90",x"14",x"E9",x"07",x"C9",x"0A",x"90", -- 0x37D0
    x"12",x"C9",x"10",x"90",x"0A",x"E9",x"20",x"C9", -- 0x37D8
    x"0A",x"90",x"08",x"C9",x"10",x"B0",x"04",x"C8", -- 0x37E0
    x"C8",x"85",x"A6",x"A5",x"F4",x"85",x"A7",x"98", -- 0x37E8
    x"48",x"A0",x"24",x"B9",x"E7",x"B8",x"99",x"52", -- 0x37F0
    x"0D",x"88",x"10",x"F7",x"A2",x"0F",x"20",x"52", -- 0x37F8
    x"0D",x"68",x"A8",x"86",x"A6",x"8A",x"10",x"14", -- 0x3800
    x"20",x"00",x"A0",x"FF",x"4E",x"6F",x"20",x"53", -- 0x3808
    x"69",x"64",x"65",x"77",x"61",x"79",x"73",x"20", -- 0x3810
    x"52",x"41",x"4D",x"00",x"20",x"62",x"82",x"18", -- 0x3818
    x"20",x"C2",x"FF",x"D0",x"03",x"4C",x"B0",x"B2", -- 0x3820
    x"20",x"FE",x"80",x"98",x"20",x"71",x"82",x"B9", -- 0x3828
    x"0E",x"0F",x"48",x"29",x"03",x"85",x"A1",x"B9", -- 0x3830
    x"0F",x"0F",x"85",x"A0",x"68",x"4A",x"4A",x"29", -- 0x3838
    x"03",x"F0",x"04",x"49",x"03",x"D0",x"16",x"B9", -- 0x3840
    x"0C",x"0F",x"D0",x"11",x"B9",x"0D",x"0F",x"30", -- 0x3848
    x"0C",x"85",x"A5",x"A2",x"05",x"C9",x"40",x"F0", -- 0x3850
    x"15",x"0A",x"CA",x"D0",x"F8",x"20",x"00",x"A0", -- 0x3858
    x"FF",x"42",x"61",x"64",x"20",x"52",x"4F",x"4D", -- 0x3860
    x"20",x"73",x"69",x"7A",x"65",x"00",x"46",x"A5", -- 0x3868
    x"A6",x"CF",x"20",x"7E",x"AA",x"18",x"A5",x"A2", -- 0x3870
    x"65",x"A0",x"85",x"A2",x"A5",x"A3",x"65",x"A1", -- 0x3878
    x"85",x"A3",x"A9",x"00",x"65",x"A4",x"85",x"A4", -- 0x3880
    x"A0",x"1C",x"B9",x"CB",x"B8",x"99",x"52",x"0D", -- 0x3888
    x"88",x"10",x"F7",x"A5",x"A6",x"8D",x"53",x"0D", -- 0x3890
    x"A5",x"A7",x"8D",x"69",x"0D",x"20",x"EC",x"A4", -- 0x3898
    x"A9",x"FF",x"8D",x"82",x"10",x"20",x"0F",x"A6", -- 0x38A0
    x"20",x"52",x"0D",x"18",x"A5",x"A2",x"69",x"02", -- 0x38A8
    x"85",x"A2",x"90",x"06",x"E6",x"A3",x"D0",x"02", -- 0x38B0
    x"E6",x"A3",x"EE",x"5E",x"0D",x"EE",x"5E",x"0D", -- 0x38B8
    x"EE",x"64",x"0D",x"EE",x"64",x"0D",x"C6",x"A5", -- 0x38C0
    x"D0",x"DB",x"60",x"A9",x"00",x"8D",x"30",x"FE", -- 0x38C8
    x"A0",x"00",x"B9",x"00",x"0E",x"99",x"00",x"80", -- 0x38D0
    x"B9",x"00",x"0F",x"99",x"00",x"81",x"88",x"D0", -- 0x38D8
    x"F1",x"A9",x"00",x"8D",x"30",x"FE",x"60",x"8E", -- 0x38E0
    x"30",x"FE",x"AD",x"FF",x"BF",x"A8",x"49",x"FF", -- 0x38E8
    x"8D",x"FF",x"BF",x"98",x"4D",x"FF",x"BF",x"8C", -- 0x38F0
    x"FF",x"BF",x"C9",x"FF",x"D0",x"04",x"C6",x"A6", -- 0x38F8
    x"30",x"03",x"CA",x"10",x"E2",x"A5",x"A7",x"8D", -- 0x3900
    x"30",x"FE",x"60",x"48",x"A5",x"CF",x"8D",x"20", -- 0x3908
    x"0D",x"68",x"60",x"A0",x"00",x"B1",x"B0",x"30", -- 0x3910
    x"07",x"29",x"03",x"85",x"CF",x"8D",x"20",x"0D", -- 0x3918
    x"A0",x"05",x"B1",x"B0",x"18",x"69",x"07",x"85", -- 0x3920
    x"BE",x"20",x"37",x"B9",x"A4",x"BE",x"B0",x"02", -- 0x3928
    x"A9",x"00",x"91",x"B0",x"A9",x"00",x"60",x"C8", -- 0x3930
    x"B1",x"B0",x"AA",x"29",x"3F",x"85",x"BF",x"C9", -- 0x3938
    x"3A",x"D0",x"2B",x"A5",x"BE",x"C9",x"09",x"D0", -- 0x3940
    x"13",x"C8",x"B1",x"B0",x"C9",x"23",x"D0",x"0C", -- 0x3948
    x"C8",x"B1",x"B0",x"29",x"20",x"F0",x"02",x"A9", -- 0x3950
    x"02",x"8D",x"20",x"0D",x"18",x"60",x"A9",x"1E", -- 0x3958
    x"38",x"60",x"A9",x"10",x"38",x"60",x"A9",x"12", -- 0x3960
    x"38",x"60",x"A9",x"FF",x"38",x"60",x"A5",x"CF", -- 0x3968
    x"6A",x"8A",x"90",x"02",x"49",x"C0",x"2A",x"90", -- 0x3970
    x"0C",x"2A",x"B0",x"E2",x"AD",x"20",x"0D",x"29", -- 0x3978
    x"02",x"09",x"01",x"D0",x"08",x"2A",x"90",x"DA", -- 0x3980
    x"AD",x"20",x"0D",x"29",x"02",x"8D",x"20",x"0D", -- 0x3988
    x"AA",x"86",x"C0",x"BD",x"10",x"0D",x"30",x"CA", -- 0x3990
    x"A5",x"BF",x"C9",x"13",x"F0",x"0B",x"C9",x"0B", -- 0x3998
    x"D0",x"BA",x"BD",x"1C",x"0D",x"C9",x"54",x"D0", -- 0x39A0
    x"BD",x"A5",x"BE",x"C9",x"0A",x"D0",x"BB",x"20", -- 0x39A8
    x"EC",x"A4",x"A9",x"00",x"85",x"C5",x"C8",x"B1", -- 0x39B0
    x"B0",x"C9",x"50",x"B0",x"A1",x"0A",x"85",x"C4", -- 0x39B8
    x"0A",x"26",x"C5",x"0A",x"26",x"C5",x"65",x"C4", -- 0x39C0
    x"85",x"C4",x"90",x"02",x"E6",x"C5",x"C8",x"B1", -- 0x39C8
    x"B0",x"C9",x"0A",x"B0",x"62",x"18",x"65",x"C4", -- 0x39D0
    x"85",x"C4",x"90",x"02",x"E6",x"C5",x"C8",x"B1", -- 0x39D8
    x"B0",x"29",x"1F",x"85",x"A5",x"F0",x"46",x"18", -- 0x39E0
    x"65",x"C4",x"AA",x"A9",x"00",x"65",x"C5",x"C9", -- 0x39E8
    x"03",x"90",x"06",x"D0",x"42",x"E0",x"21",x"B0", -- 0x39F0
    x"3E",x"A6",x"C0",x"BD",x"10",x"0D",x"6A",x"BD", -- 0x39F8
    x"0C",x"0D",x"20",x"87",x"AA",x"18",x"A5",x"A2", -- 0x3A00
    x"65",x"C4",x"85",x"A2",x"A5",x"A3",x"65",x"C5", -- 0x3A08
    x"85",x"A3",x"90",x"02",x"E6",x"A4",x"A0",x"00", -- 0x3A10
    x"84",x"A7",x"C8",x"B1",x"B0",x"85",x"A0",x"C8", -- 0x3A18
    x"B1",x"B0",x"85",x"A1",x"A5",x"BF",x"C9",x"13", -- 0x3A20
    x"F0",x"05",x"20",x"AB",x"AB",x"18",x"60",x"20", -- 0x3A28
    x"42",x"A6",x"20",x"CD",x"A0",x"18",x"60",x"A9", -- 0x3A30
    x"1E",x"38",x"60",x"54",x"45",x"53",x"53",x"20", -- 0x3A38
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3A40
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3A48
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3A50
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3A58
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3A60
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3A68
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3A70
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3A78
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3A80
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3A88
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3A90
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3A98
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3AA0
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3AA8
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3AB0
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3AB8
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3AC0
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3AC8
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3AD0
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3AD8
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3AE0
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3AE8
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3AF0
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3AF8
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3B00
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3B08
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3B10
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3B18
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3B20
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3B28
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3B30
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3B38
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3B40
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3B48
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3B50
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3B58
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3B60
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3B68
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3B70
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3B78
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3B80
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3B88
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3B90
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3B98
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3BA0
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3BA8
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3BB0
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3BB8
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3BC0
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3BC8
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3BD0
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3BD8
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3BE0
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3BE8
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3BF0
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3BF8
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3C00
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3C08
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3C10
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3C18
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3C20
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3C28
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3C30
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3C38
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3C40
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3C48
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3C50
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3C58
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3C60
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3C68
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3C70
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3C78
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3C80
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3C88
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3C90
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3C98
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3CA0
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3CA8
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3CB0
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3CB8
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3CC0
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3CC8
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3CD0
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3CD8
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3CE0
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3CE8
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3CF0
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3CF8
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3D00
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3D08
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3D10
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3D18
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3D20
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3D28
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3D30
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3D38
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3D40
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3D48
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3D50
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3D58
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3D60
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3D68
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3D70
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3D78
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3D80
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3D88
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3D90
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3D98
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3DA0
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3DA8
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3DB0
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3DB8
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3DC0
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3DC8
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3DD0
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3DD8
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3DE0
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3DE8
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3DF0
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3DF8
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3E00
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3E08
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3E10
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3E18
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3E20
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3E28
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3E30
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3E38
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3E40
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3E48
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3E50
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3E58
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3E60
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3E68
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3E70
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3E78
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3E80
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3E88
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3E90
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3E98
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3EA0
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3EA8
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3EB0
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3EB8
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3EC0
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3EC8
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3ED0
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3ED8
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3EE0
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3EE8
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3EF0
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3EF8
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3F00
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3F08
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3F10
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3F18
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3F20
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3F28
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3F30
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3F38
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3F40
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3F48
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3F50
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3F58
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3F60
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3F68
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3F70
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3F78
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3F80
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3F88
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3F90
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3F98
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3FA0
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3FA8
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3FB0
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3FB8
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3FC0
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3FC8
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45", -- 0x3FD0
    x"53",x"53",x"20",x"54",x"45",x"53",x"53",x"20", -- 0x3FD8
    x"54",x"45",x"53",x"53",x"20",x"54",x"45",x"53", -- 0x3FE0
    x"53",x"20",x"54",x"45",x"53",x"53",x"20",x"54", -- 0x3FE8
    x"45",x"53",x"53",x"20",x"54",x"45",x"53",x"53", -- 0x3FF0
    x"20",x"54",x"45",x"53",x"53",x"20",x"54",x"45"  -- 0x3FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
     DATA <= ROM(to_integer(unsigned(ADDR)));
  end process;
end RTL;
