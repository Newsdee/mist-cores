-- generated with romgen by MikeJ
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity BBC_OS12_ROM is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of BBC_OS12_ROM is


  type ROM_ARRAY is array(0 to 16383) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0000
    x"18",x"18",x"18",x"18",x"18",x"00",x"18",x"00", -- 0x0008
    x"6C",x"6C",x"6C",x"00",x"00",x"00",x"00",x"00", -- 0x0010
    x"36",x"36",x"7F",x"36",x"7F",x"36",x"36",x"00", -- 0x0018
    x"0C",x"3F",x"68",x"3E",x"0B",x"7E",x"18",x"00", -- 0x0020
    x"60",x"66",x"0C",x"18",x"30",x"66",x"06",x"00", -- 0x0028
    x"38",x"6C",x"6C",x"38",x"6D",x"66",x"3B",x"00", -- 0x0030
    x"0C",x"18",x"30",x"00",x"00",x"00",x"00",x"00", -- 0x0038
    x"0C",x"18",x"30",x"30",x"30",x"18",x"0C",x"00", -- 0x0040
    x"30",x"18",x"0C",x"0C",x"0C",x"18",x"30",x"00", -- 0x0048
    x"00",x"18",x"7E",x"3C",x"7E",x"18",x"00",x"00", -- 0x0050
    x"00",x"18",x"18",x"7E",x"18",x"18",x"00",x"00", -- 0x0058
    x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"30", -- 0x0060
    x"00",x"00",x"00",x"7E",x"00",x"00",x"00",x"00", -- 0x0068
    x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00", -- 0x0070
    x"00",x"06",x"0C",x"18",x"30",x"60",x"00",x"00", -- 0x0078
    x"3C",x"66",x"6E",x"7E",x"76",x"66",x"3C",x"00", -- 0x0080
    x"18",x"38",x"18",x"18",x"18",x"18",x"7E",x"00", -- 0x0088
    x"3C",x"66",x"06",x"0C",x"18",x"30",x"7E",x"00", -- 0x0090
    x"3C",x"66",x"06",x"1C",x"06",x"66",x"3C",x"00", -- 0x0098
    x"0C",x"1C",x"3C",x"6C",x"7E",x"0C",x"0C",x"00", -- 0x00A0
    x"7E",x"60",x"7C",x"06",x"06",x"66",x"3C",x"00", -- 0x00A8
    x"1C",x"30",x"60",x"7C",x"66",x"66",x"3C",x"00", -- 0x00B0
    x"7E",x"06",x"0C",x"18",x"30",x"30",x"30",x"00", -- 0x00B8
    x"3C",x"66",x"66",x"3C",x"66",x"66",x"3C",x"00", -- 0x00C0
    x"3C",x"66",x"66",x"3E",x"06",x"0C",x"38",x"00", -- 0x00C8
    x"00",x"00",x"18",x"18",x"00",x"18",x"18",x"00", -- 0x00D0
    x"00",x"00",x"18",x"18",x"00",x"18",x"18",x"30", -- 0x00D8
    x"0C",x"18",x"30",x"60",x"30",x"18",x"0C",x"00", -- 0x00E0
    x"00",x"00",x"7E",x"00",x"7E",x"00",x"00",x"00", -- 0x00E8
    x"30",x"18",x"0C",x"06",x"0C",x"18",x"30",x"00", -- 0x00F0
    x"3C",x"66",x"0C",x"18",x"18",x"00",x"18",x"00", -- 0x00F8
    x"3C",x"66",x"6E",x"6A",x"6E",x"60",x"3C",x"00", -- 0x0100
    x"3C",x"66",x"66",x"7E",x"66",x"66",x"66",x"00", -- 0x0108
    x"7C",x"66",x"66",x"7C",x"66",x"66",x"7C",x"00", -- 0x0110
    x"3C",x"66",x"60",x"60",x"60",x"66",x"3C",x"00", -- 0x0118
    x"78",x"6C",x"66",x"66",x"66",x"6C",x"78",x"00", -- 0x0120
    x"7E",x"60",x"60",x"7C",x"60",x"60",x"7E",x"00", -- 0x0128
    x"7E",x"60",x"60",x"7C",x"60",x"60",x"60",x"00", -- 0x0130
    x"3C",x"66",x"60",x"6E",x"66",x"66",x"3C",x"00", -- 0x0138
    x"66",x"66",x"66",x"7E",x"66",x"66",x"66",x"00", -- 0x0140
    x"7E",x"18",x"18",x"18",x"18",x"18",x"7E",x"00", -- 0x0148
    x"3E",x"0C",x"0C",x"0C",x"0C",x"6C",x"38",x"00", -- 0x0150
    x"66",x"6C",x"78",x"70",x"78",x"6C",x"66",x"00", -- 0x0158
    x"60",x"60",x"60",x"60",x"60",x"60",x"7E",x"00", -- 0x0160
    x"63",x"77",x"7F",x"6B",x"6B",x"63",x"63",x"00", -- 0x0168
    x"66",x"66",x"76",x"7E",x"6E",x"66",x"66",x"00", -- 0x0170
    x"3C",x"66",x"66",x"66",x"66",x"66",x"3C",x"00", -- 0x0178
    x"7C",x"66",x"66",x"7C",x"60",x"60",x"60",x"00", -- 0x0180
    x"3C",x"66",x"66",x"66",x"6A",x"6C",x"36",x"00", -- 0x0188
    x"7C",x"66",x"66",x"7C",x"6C",x"66",x"66",x"00", -- 0x0190
    x"3C",x"66",x"60",x"3C",x"06",x"66",x"3C",x"00", -- 0x0198
    x"7E",x"18",x"18",x"18",x"18",x"18",x"18",x"00", -- 0x01A0
    x"66",x"66",x"66",x"66",x"66",x"66",x"3C",x"00", -- 0x01A8
    x"66",x"66",x"66",x"66",x"66",x"3C",x"18",x"00", -- 0x01B0
    x"63",x"63",x"6B",x"6B",x"7F",x"77",x"63",x"00", -- 0x01B8
    x"66",x"66",x"3C",x"18",x"3C",x"66",x"66",x"00", -- 0x01C0
    x"66",x"66",x"66",x"3C",x"18",x"18",x"18",x"00", -- 0x01C8
    x"7E",x"06",x"0C",x"18",x"30",x"60",x"7E",x"00", -- 0x01D0
    x"7C",x"60",x"60",x"60",x"60",x"60",x"7C",x"00", -- 0x01D8
    x"00",x"60",x"30",x"18",x"0C",x"06",x"00",x"00", -- 0x01E0
    x"3E",x"06",x"06",x"06",x"06",x"06",x"3E",x"00", -- 0x01E8
    x"18",x"3C",x"66",x"42",x"00",x"00",x"00",x"00", -- 0x01F0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF", -- 0x01F8
    x"1C",x"36",x"30",x"7C",x"30",x"30",x"7E",x"00", -- 0x0200
    x"00",x"00",x"3C",x"06",x"3E",x"66",x"3E",x"00", -- 0x0208
    x"60",x"60",x"7C",x"66",x"66",x"66",x"7C",x"00", -- 0x0210
    x"00",x"00",x"3C",x"66",x"60",x"66",x"3C",x"00", -- 0x0218
    x"06",x"06",x"3E",x"66",x"66",x"66",x"3E",x"00", -- 0x0220
    x"00",x"00",x"3C",x"66",x"7E",x"60",x"3C",x"00", -- 0x0228
    x"1C",x"30",x"30",x"7C",x"30",x"30",x"30",x"00", -- 0x0230
    x"00",x"00",x"3E",x"66",x"66",x"3E",x"06",x"3C", -- 0x0238
    x"60",x"60",x"7C",x"66",x"66",x"66",x"66",x"00", -- 0x0240
    x"18",x"00",x"38",x"18",x"18",x"18",x"3C",x"00", -- 0x0248
    x"18",x"00",x"38",x"18",x"18",x"18",x"18",x"70", -- 0x0250
    x"60",x"60",x"66",x"6C",x"78",x"6C",x"66",x"00", -- 0x0258
    x"38",x"18",x"18",x"18",x"18",x"18",x"3C",x"00", -- 0x0260
    x"00",x"00",x"36",x"7F",x"6B",x"6B",x"63",x"00", -- 0x0268
    x"00",x"00",x"7C",x"66",x"66",x"66",x"66",x"00", -- 0x0270
    x"00",x"00",x"3C",x"66",x"66",x"66",x"3C",x"00", -- 0x0278
    x"00",x"00",x"7C",x"66",x"66",x"7C",x"60",x"60", -- 0x0280
    x"00",x"00",x"3E",x"66",x"66",x"3E",x"06",x"07", -- 0x0288
    x"00",x"00",x"6C",x"76",x"60",x"60",x"60",x"00", -- 0x0290
    x"00",x"00",x"3E",x"60",x"3C",x"06",x"7C",x"00", -- 0x0298
    x"30",x"30",x"7C",x"30",x"30",x"30",x"1C",x"00", -- 0x02A0
    x"00",x"00",x"66",x"66",x"66",x"66",x"3E",x"00", -- 0x02A8
    x"00",x"00",x"66",x"66",x"66",x"3C",x"18",x"00", -- 0x02B0
    x"00",x"00",x"63",x"6B",x"6B",x"7F",x"36",x"00", -- 0x02B8
    x"00",x"00",x"66",x"3C",x"18",x"3C",x"66",x"00", -- 0x02C0
    x"00",x"00",x"66",x"66",x"66",x"3E",x"06",x"3C", -- 0x02C8
    x"00",x"00",x"7E",x"0C",x"18",x"30",x"7E",x"00", -- 0x02D0
    x"0C",x"18",x"18",x"70",x"18",x"18",x"0C",x"00", -- 0x02D8
    x"18",x"18",x"18",x"00",x"18",x"18",x"18",x"00", -- 0x02E0
    x"30",x"18",x"18",x"0E",x"18",x"18",x"30",x"00", -- 0x02E8
    x"31",x"6B",x"46",x"00",x"00",x"00",x"00",x"00", -- 0x02F0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02F8
    x"4C",x"1D",x"CB",x"0D",x"42",x"42",x"43",x"20", -- 0x0300
    x"43",x"6F",x"6D",x"70",x"75",x"74",x"65",x"72", -- 0x0308
    x"20",x"00",x"31",x"36",x"4B",x"07",x"00",x"33", -- 0x0310
    x"32",x"4B",x"07",x"00",x"08",x"0D",x"0D",x"00", -- 0x0318
    x"11",x"22",x"33",x"44",x"55",x"66",x"77",x"88", -- 0x0320
    x"99",x"AA",x"BB",x"CC",x"DD",x"EE",x"FF",x"00", -- 0x0328
    x"55",x"AA",x"FF",x"11",x"3B",x"96",x"A1",x"AD", -- 0x0330
    x"B9",x"11",x"6F",x"C5",x"64",x"F0",x"5B",x"59", -- 0x0338
    x"AF",x"8D",x"A6",x"C0",x"F9",x"FD",x"92",x"39", -- 0x0340
    x"9B",x"EB",x"F1",x"39",x"8C",x"BD",x"11",x"FA", -- 0x0348
    x"A2",x"79",x"87",x"AC",x"C5",x"2F",x"C5",x"C5", -- 0x0350
    x"C5",x"C5",x"C5",x"E8",x"C5",x"C6",x"C6",x"C6", -- 0x0358
    x"C7",x"C7",x"C5",x"C5",x"C7",x"4F",x"4E",x"5B", -- 0x0360
    x"C8",x"C5",x"5F",x"57",x"78",x"6B",x"C9",x"C5", -- 0x0368
    x"3C",x"7C",x"C7",x"4E",x"CA",x"00",x"00",x"02", -- 0x0370
    x"80",x"05",x"00",x"07",x"80",x"0A",x"00",x"0C", -- 0x0378
    x"80",x"0F",x"00",x"11",x"80",x"14",x"00",x"16", -- 0x0380
    x"80",x"19",x"00",x"1B",x"80",x"1E",x"00",x"20", -- 0x0388
    x"80",x"23",x"00",x"25",x"80",x"28",x"00",x"2A", -- 0x0390
    x"80",x"2D",x"00",x"2F",x"80",x"32",x"00",x"34", -- 0x0398
    x"80",x"37",x"00",x"39",x"80",x"3C",x"00",x"3E", -- 0x03A0
    x"80",x"41",x"00",x"43",x"80",x"46",x"00",x"48", -- 0x03A8
    x"80",x"4B",x"00",x"4D",x"80",x"00",x"00",x"00", -- 0x03B0
    x"28",x"00",x"50",x"00",x"78",x"00",x"A0",x"00", -- 0x03B8
    x"C8",x"00",x"F0",x"01",x"18",x"01",x"40",x"01", -- 0x03C0
    x"68",x"01",x"90",x"01",x"B8",x"01",x"E0",x"02", -- 0x03C8
    x"08",x"02",x"30",x"02",x"58",x"02",x"80",x"02", -- 0x03D0
    x"A8",x"02",x"D0",x"02",x"F8",x"03",x"20",x"03", -- 0x03D8
    x"48",x"03",x"70",x"03",x"98",x"03",x"C0",x"1F", -- 0x03E0
    x"1F",x"1F",x"18",x"1F",x"1F",x"18",x"18",x"4F", -- 0x03E8
    x"27",x"13",x"4F",x"27",x"13",x"27",x"27",x"9C", -- 0x03F0
    x"D8",x"F4",x"9C",x"88",x"C4",x"88",x"4B",x"08", -- 0x03F8
    x"10",x"20",x"08",x"08",x"10",x"08",x"01",x"AA", -- 0x0400
    x"55",x"88",x"44",x"22",x"11",x"80",x"40",x"20", -- 0x0408
    x"10",x"08",x"04",x"02",x"01",x"03",x"0F",x"01", -- 0x0410
    x"01",x"03",x"01",x"00",x"FF",x"00",x"00",x"FF", -- 0x0418
    x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"00",x"0F", -- 0x0420
    x"F0",x"FF",x"00",x"03",x"0C",x"0F",x"30",x"33", -- 0x0428
    x"3C",x"3F",x"C0",x"C3",x"CC",x"CF",x"F0",x"F3", -- 0x0430
    x"FC",x"FF",x"07",x"03",x"01",x"00",x"07",x"03", -- 0x0438
    x"00",x"00",x"00",x"01",x"02",x"02",x"03",x"04", -- 0x0440
    x"00",x"06",x"02",x"0D",x"05",x"0D",x"05",x"04", -- 0x0448
    x"04",x"0C",x"0C",x"04",x"02",x"32",x"7A",x"92", -- 0x0450
    x"E6",x"50",x"40",x"28",x"20",x"04",x"30",x"40", -- 0x0458
    x"58",x"60",x"7C",x"28",x"40",x"80",x"B5",x"75", -- 0x0460
    x"75",x"0B",x"17",x"23",x"2F",x"3B",x"7F",x"50", -- 0x0468
    x"62",x"28",x"26",x"00",x"20",x"22",x"01",x"07", -- 0x0470
    x"67",x"08",x"7F",x"50",x"62",x"28",x"1E",x"02", -- 0x0478
    x"19",x"1B",x"01",x"09",x"67",x"09",x"3F",x"28", -- 0x0480
    x"31",x"24",x"26",x"00",x"20",x"22",x"01",x"07", -- 0x0488
    x"67",x"08",x"3F",x"28",x"31",x"24",x"1E",x"02", -- 0x0490
    x"19",x"1B",x"01",x"09",x"67",x"09",x"3F",x"28", -- 0x0498
    x"33",x"24",x"1E",x"02",x"19",x"1B",x"93",x"12", -- 0x04A0
    x"72",x"13",x"86",x"D3",x"7E",x"D3",x"6A",x"74", -- 0x04A8
    x"42",x"4B",x"D3",x"D3",x"D3",x"D3",x"23",x"5F", -- 0x04B0
    x"60",x"23",x"04",x"05",x"06",x"00",x"01",x"02", -- 0x04B8
    x"AE",x"6A",x"02",x"D0",x"4D",x"24",x"D0",x"50", -- 0x04C0
    x"0F",x"20",x"68",x"C5",x"20",x"6A",x"CD",x"30", -- 0x04C8
    x"07",x"C9",x"0D",x"D0",x"03",x"20",x"18",x"D9", -- 0x04D0
    x"C9",x"7F",x"F0",x"11",x"C9",x"20",x"90",x"0F", -- 0x04D8
    x"24",x"D0",x"30",x"06",x"20",x"B7",x"CF",x"20", -- 0x04E0
    x"64",x"C6",x"4C",x"5E",x"C5",x"A9",x"20",x"A8", -- 0x04E8
    x"B9",x"33",x"C3",x"8D",x"5D",x"03",x"B9",x"54", -- 0x04F0
    x"C3",x"30",x"4A",x"AA",x"09",x"F0",x"8D",x"6A", -- 0x04F8
    x"02",x"8A",x"4A",x"4A",x"4A",x"4A",x"18",x"69", -- 0x0500
    x"C3",x"8D",x"5E",x"03",x"24",x"D0",x"70",x"1F", -- 0x0508
    x"18",x"60",x"9D",x"24",x"02",x"E8",x"8E",x"6A", -- 0x0510
    x"02",x"D0",x"17",x"24",x"D0",x"30",x"15",x"70", -- 0x0518
    x"05",x"20",x"F5",x"CC",x"18",x"60",x"20",x"68", -- 0x0520
    x"C5",x"20",x"6A",x"CD",x"20",x"F5",x"CC",x"20", -- 0x0528
    x"65",x"C5",x"18",x"60",x"AC",x"5E",x"03",x"C0", -- 0x0530
    x"C5",x"D0",x"F7",x"AA",x"A5",x"D0",x"4A",x"90", -- 0x0538
    x"D0",x"8A",x"4C",x"1E",x"E1",x"8D",x"5E",x"03", -- 0x0540
    x"98",x"C9",x"08",x"90",x"06",x"49",x"FF",x"C9", -- 0x0548
    x"F2",x"49",x"FF",x"24",x"D0",x"30",x"29",x"08", -- 0x0550
    x"20",x"F5",x"CC",x"28",x"90",x"03",x"A5",x"D0", -- 0x0558
    x"4A",x"24",x"D0",x"50",x"AC",x"20",x"7A",x"CD", -- 0x0560
    x"08",x"48",x"A2",x"18",x"A0",x"64",x"20",x"DE", -- 0x0568
    x"CD",x"20",x"06",x"CF",x"20",x"02",x"CA",x"A5", -- 0x0570
    x"D0",x"49",x"02",x"85",x"D0",x"68",x"28",x"60", -- 0x0578
    x"49",x"06",x"D0",x"08",x"A9",x"7F",x"90",x"20", -- 0x0580
    x"A5",x"D0",x"29",x"20",x"60",x"A0",x"00",x"8C", -- 0x0588
    x"69",x"02",x"A9",x"04",x"D0",x"07",x"20",x"A2", -- 0x0590
    x"E1",x"A9",x"94",x"49",x"95",x"05",x"D0",x"D0", -- 0x0598
    x"09",x"20",x"A2",x"E1",x"A9",x"0A",x"49",x"F4", -- 0x05A0
    x"25",x"D0",x"85",x"D0",x"60",x"AD",x"61",x"03", -- 0x05A8
    x"F0",x"FA",x"20",x"51",x"C9",x"A9",x"DF",x"D0", -- 0x05B0
    x"EF",x"AD",x"61",x"03",x"F0",x"EE",x"A9",x"20", -- 0x05B8
    x"20",x"54",x"C9",x"D0",x"D8",x"20",x"88",x"C5", -- 0x05C0
    x"D0",x"55",x"CE",x"18",x"03",x"AE",x"18",x"03", -- 0x05C8
    x"EC",x"08",x"03",x"30",x"19",x"AD",x"4A",x"03", -- 0x05D0
    x"38",x"ED",x"4F",x"03",x"AA",x"AD",x"4B",x"03", -- 0x05D8
    x"E9",x"00",x"CD",x"4E",x"03",x"B0",x"03",x"6D", -- 0x05E0
    x"54",x"03",x"A8",x"4C",x"F6",x"C9",x"AD",x"0A", -- 0x05E8
    x"03",x"8D",x"18",x"03",x"CE",x"69",x"02",x"10", -- 0x05F0
    x"03",x"EE",x"69",x"02",x"AE",x"19",x"03",x"EC", -- 0x05F8
    x"0B",x"03",x"F0",x"06",x"CE",x"19",x"03",x"4C", -- 0x0600
    x"AF",x"C6",x"18",x"20",x"3F",x"CD",x"A9",x"08", -- 0x0608
    x"24",x"D0",x"D0",x"05",x"20",x"94",x"C9",x"D0", -- 0x0610
    x"03",x"20",x"A4",x"CD",x"4C",x"AC",x"C6",x"A2", -- 0x0618
    x"00",x"86",x"DB",x"20",x"0D",x"D1",x"A6",x"DB", -- 0x0620
    x"38",x"BD",x"24",x"03",x"E9",x"08",x"9D",x"24", -- 0x0628
    x"03",x"B0",x"03",x"DE",x"25",x"03",x"A5",x"DA", -- 0x0630
    x"D0",x"1E",x"20",x"0D",x"D1",x"F0",x"19",x"A6", -- 0x0638
    x"DB",x"BD",x"04",x"03",x"E0",x"01",x"B0",x"02", -- 0x0640
    x"E9",x"06",x"9D",x"24",x"03",x"BD",x"05",x"03", -- 0x0648
    x"E9",x"00",x"9D",x"25",x"03",x"8A",x"F0",x"08", -- 0x0650
    x"4C",x"B8",x"D1",x"20",x"88",x"C5",x"F0",x"94", -- 0x0658
    x"A2",x"02",x"D0",x"52",x"A5",x"D0",x"29",x"20", -- 0x0660
    x"D0",x"4A",x"AE",x"18",x"03",x"EC",x"0A",x"03", -- 0x0668
    x"B0",x"12",x"EE",x"18",x"03",x"AD",x"4A",x"03", -- 0x0670
    x"6D",x"4F",x"03",x"AA",x"AD",x"4B",x"03",x"69", -- 0x0678
    x"00",x"4C",x"F6",x"C9",x"AD",x"08",x"03",x"8D", -- 0x0680
    x"18",x"03",x"18",x"20",x"E3",x"CA",x"AE",x"19", -- 0x0688
    x"03",x"EC",x"09",x"03",x"B0",x"05",x"EE",x"19", -- 0x0690
    x"03",x"90",x"14",x"20",x"3F",x"CD",x"A9",x"08", -- 0x0698
    x"24",x"D0",x"D0",x"05",x"20",x"A4",x"C9",x"D0", -- 0x06A0
    x"03",x"20",x"FF",x"CD",x"20",x"AC",x"CE",x"20", -- 0x06A8
    x"06",x"CF",x"90",x"7E",x"A2",x"00",x"86",x"DB", -- 0x06B0
    x"20",x"0D",x"D1",x"A6",x"DB",x"18",x"BD",x"24", -- 0x06B8
    x"03",x"69",x"08",x"9D",x"24",x"03",x"90",x"03", -- 0x06C0
    x"FE",x"25",x"03",x"A5",x"DA",x"D0",x"89",x"20", -- 0x06C8
    x"0D",x"D1",x"F0",x"84",x"A6",x"DB",x"BD",x"00", -- 0x06D0
    x"03",x"E0",x"01",x"90",x"02",x"69",x"06",x"9D", -- 0x06D8
    x"24",x"03",x"BD",x"01",x"03",x"69",x"00",x"9D", -- 0x06E0
    x"25",x"03",x"8A",x"F0",x"08",x"4C",x"B8",x"D1", -- 0x06E8
    x"20",x"88",x"C5",x"F0",x"95",x"A2",x"02",x"4C", -- 0x06F0
    x"21",x"C6",x"AE",x"55",x"03",x"AD",x"21",x"03", -- 0x06F8
    x"CD",x"23",x"03",x"90",x"53",x"DD",x"E7",x"C3", -- 0x0700
    x"F0",x"02",x"B0",x"4C",x"AD",x"22",x"03",x"A8", -- 0x0708
    x"DD",x"EF",x"C3",x"F0",x"02",x"B0",x"41",x"38", -- 0x0710
    x"ED",x"20",x"03",x"30",x"3B",x"A8",x"20",x"88", -- 0x0718
    x"CA",x"A9",x"08",x"20",x"9D",x"C5",x"A2",x"20", -- 0x0720
    x"A0",x"08",x"20",x"8A",x"D4",x"20",x"E8",x"CE", -- 0x0728
    x"B0",x"47",x"4C",x"02",x"CA",x"A0",x"03",x"B1", -- 0x0730
    x"F0",x"99",x"28",x"03",x"88",x"10",x"F8",x"A9", -- 0x0738
    x"28",x"20",x"39",x"D8",x"A0",x"04",x"D0",x"08", -- 0x0740
    x"2D",x"60",x"03",x"AA",x"BD",x"6F",x"03",x"C8", -- 0x0748
    x"91",x"F0",x"A9",x"00",x"C0",x"04",x"D0",x"F7", -- 0x0750
    x"60",x"20",x"88",x"C5",x"D0",x"5F",x"A5",x"D0", -- 0x0758
    x"29",x"08",x"D0",x"03",x"4C",x"C1",x"CB",x"AE", -- 0x0760
    x"0B",x"03",x"8E",x"19",x"03",x"20",x"AC",x"CE", -- 0x0768
    x"AE",x"19",x"03",x"EC",x"09",x"03",x"E8",x"90", -- 0x0770
    x"F1",x"20",x"88",x"C5",x"F0",x"03",x"4C",x"A6", -- 0x0778
    x"CF",x"8D",x"23",x"03",x"8D",x"22",x"03",x"20", -- 0x0780
    x"88",x"C5",x"D0",x"CC",x"20",x"A8",x"C7",x"18", -- 0x0788
    x"AD",x"22",x"03",x"6D",x"08",x"03",x"8D",x"18", -- 0x0790
    x"03",x"AD",x"23",x"03",x"18",x"6D",x"0B",x"03", -- 0x0798
    x"8D",x"19",x"03",x"20",x"E8",x"CE",x"90",x"8A", -- 0x07A0
    x"A2",x"18",x"A0",x"28",x"4C",x"DE",x"CD",x"20", -- 0x07A8
    x"88",x"C5",x"F0",x"03",x"4C",x"AD",x"CF",x"20", -- 0x07B0
    x"6E",x"CE",x"4C",x"AF",x"C6",x"20",x"A6",x"CF", -- 0x07B8
    x"AD",x"61",x"03",x"F0",x"33",x"AE",x"5A",x"03", -- 0x07C0
    x"AC",x"5C",x"03",x"20",x"B3",x"D0",x"A2",x"00", -- 0x07C8
    x"A0",x"28",x"20",x"7C",x"D4",x"38",x"AD",x"06", -- 0x07D0
    x"03",x"ED",x"02",x"03",x"A8",x"C8",x"8C",x"30", -- 0x07D8
    x"03",x"A2",x"2C",x"A0",x"28",x"20",x"A6",x"D6", -- 0x07E0
    x"AD",x"2E",x"03",x"D0",x"03",x"CE",x"2F",x"03", -- 0x07E8
    x"CE",x"2E",x"03",x"CE",x"30",x"03",x"D0",x"E9", -- 0x07F0
    x"60",x"A0",x"00",x"F0",x"02",x"A0",x"02",x"AD", -- 0x07F8
    x"23",x"03",x"10",x"01",x"C8",x"2D",x"60",x"03", -- 0x0800
    x"85",x"DA",x"AD",x"60",x"03",x"F0",x"1C",x"29", -- 0x0808
    x"07",x"18",x"65",x"DA",x"AA",x"BD",x"23",x"C4", -- 0x0810
    x"99",x"57",x"03",x"C0",x"02",x"B0",x"0D",x"AD", -- 0x0818
    x"57",x"03",x"49",x"FF",x"85",x"D3",x"4D",x"58", -- 0x0820
    x"03",x"85",x"D2",x"60",x"AD",x"22",x"03",x"99", -- 0x0828
    x"59",x"03",x"60",x"A9",x"20",x"8D",x"58",x"03", -- 0x0830
    x"60",x"A2",x"05",x"A9",x"00",x"9D",x"57",x"03", -- 0x0838
    x"CA",x"10",x"FA",x"AE",x"60",x"03",x"F0",x"EB", -- 0x0840
    x"A9",x"FF",x"E0",x"0F",x"D0",x"02",x"A9",x"3F", -- 0x0848
    x"8D",x"57",x"03",x"8D",x"59",x"03",x"49",x"FF", -- 0x0850
    x"85",x"D2",x"85",x"D3",x"8E",x"1F",x"03",x"E0", -- 0x0858
    x"03",x"F0",x"11",x"90",x"20",x"8E",x"20",x"03", -- 0x0860
    x"20",x"92",x"C8",x"CE",x"20",x"03",x"CE",x"1F", -- 0x0868
    x"03",x"10",x"F5",x"60",x"A2",x"07",x"8E",x"20", -- 0x0870
    x"03",x"20",x"92",x"C8",x"4E",x"20",x"03",x"CE", -- 0x0878
    x"1F",x"03",x"10",x"F5",x"60",x"A2",x"07",x"20", -- 0x0880
    x"8F",x"C8",x"A2",x"00",x"8E",x"1F",x"03",x"8E", -- 0x0888
    x"20",x"03",x"08",x"78",x"AD",x"1F",x"03",x"2D", -- 0x0890
    x"60",x"03",x"AA",x"AD",x"20",x"03",x"29",x"0F", -- 0x0898
    x"9D",x"6F",x"03",x"A8",x"AD",x"60",x"03",x"85", -- 0x08A0
    x"FA",x"C9",x"03",x"08",x"8A",x"6A",x"66",x"FA", -- 0x08A8
    x"B0",x"FB",x"06",x"FA",x"98",x"05",x"FA",x"AA", -- 0x08B0
    x"A0",x"00",x"28",x"08",x"D0",x"0E",x"29",x"60", -- 0x08B8
    x"F0",x"09",x"C9",x"60",x"F0",x"05",x"8A",x"49", -- 0x08C0
    x"60",x"D0",x"01",x"8A",x"20",x"11",x"EA",x"98", -- 0x08C8
    x"38",x"6D",x"60",x"03",x"A8",x"8A",x"69",x"10", -- 0x08D0
    x"AA",x"C0",x"10",x"90",x"DD",x"28",x"28",x"60", -- 0x08D8
    x"08",x"2D",x"60",x"03",x"AA",x"C8",x"B1",x"F0", -- 0x08E0
    x"4C",x"9E",x"C8",x"AD",x"23",x"03",x"4C",x"33", -- 0x08E8
    x"CB",x"AD",x"1B",x"03",x"C9",x"20",x"90",x"47", -- 0x08F0
    x"48",x"4A",x"4A",x"4A",x"4A",x"4A",x"AA",x"BD", -- 0x08F8
    x"0D",x"C4",x"2C",x"67",x"03",x"D0",x"20",x"0D", -- 0x0900
    x"67",x"03",x"8D",x"67",x"03",x"8A",x"29",x"03", -- 0x0908
    x"18",x"69",x"BF",x"85",x"DF",x"BD",x"67",x"03", -- 0x0910
    x"85",x"DD",x"A0",x"00",x"84",x"DC",x"84",x"DE", -- 0x0918
    x"B1",x"DE",x"91",x"DC",x"88",x"D0",x"F9",x"68", -- 0x0920
    x"20",x"3E",x"D0",x"A0",x"07",x"B9",x"1C",x"03", -- 0x0928
    x"91",x"DE",x"88",x"10",x"F8",x"60",x"68",x"60", -- 0x0930
    x"AD",x"1F",x"03",x"18",x"6C",x"26",x"02",x"C9", -- 0x0938
    x"01",x"90",x"15",x"D0",x"F7",x"20",x"88",x"C5", -- 0x0940
    x"D0",x"ED",x"A9",x"20",x"AC",x"1C",x"03",x"F0", -- 0x0948
    x"03",x"AD",x"5F",x"03",x"A0",x"0A",x"D0",x"2D", -- 0x0950
    x"AD",x"1D",x"03",x"AC",x"1C",x"03",x"C0",x"07", -- 0x0958
    x"90",x"23",x"D0",x"03",x"6D",x"90",x"02",x"C0", -- 0x0960
    x"08",x"D0",x"07",x"09",x"00",x"30",x"03",x"4D", -- 0x0968
    x"91",x"02",x"C0",x"0A",x"D0",x"0F",x"8D",x"5F", -- 0x0970
    x"03",x"A8",x"A5",x"D0",x"29",x"20",x"08",x"98", -- 0x0978
    x"A0",x"0A",x"28",x"D0",x"06",x"8C",x"00",x"FE", -- 0x0980
    x"8D",x"01",x"FE",x"60",x"AE",x"61",x"03",x"F0", -- 0x0988
    x"A7",x"4C",x"60",x"D0",x"AE",x"50",x"03",x"AD", -- 0x0990
    x"51",x"03",x"20",x"F8",x"CC",x"B0",x"14",x"6D", -- 0x0998
    x"54",x"03",x"90",x"0F",x"AE",x"50",x"03",x"AD", -- 0x09A0
    x"51",x"03",x"20",x"D4",x"CA",x"10",x"04",x"38", -- 0x09A8
    x"ED",x"54",x"03",x"8D",x"51",x"03",x"8E",x"50", -- 0x09B0
    x"03",x"A0",x"0C",x"D0",x"51",x"A9",x"00",x"A2", -- 0x09B8
    x"2C",x"9D",x"00",x"03",x"CA",x"10",x"FA",x"AE", -- 0x09C0
    x"55",x"03",x"BC",x"EF",x"C3",x"8C",x"0A",x"03", -- 0x09C8
    x"20",x"88",x"CA",x"BC",x"E7",x"C3",x"8C",x"09", -- 0x09D0
    x"03",x"A0",x"03",x"8C",x"23",x"03",x"C8",x"8C", -- 0x09D8
    x"21",x"03",x"CE",x"22",x"03",x"CE",x"20",x"03", -- 0x09E0
    x"20",x"39",x"CA",x"A9",x"F7",x"20",x"A8",x"C5", -- 0x09E8
    x"AE",x"50",x"03",x"AD",x"51",x"03",x"8E",x"4A", -- 0x09F0
    x"03",x"8D",x"4B",x"03",x"10",x"04",x"38",x"ED", -- 0x09F8
    x"54",x"03",x"86",x"D8",x"85",x"D9",x"AE",x"4A", -- 0x0A00
    x"03",x"AD",x"4B",x"03",x"A0",x"0E",x"48",x"AD", -- 0x0A08
    x"55",x"03",x"C9",x"07",x"68",x"B0",x"10",x"86", -- 0x0A10
    x"DA",x"4A",x"66",x"DA",x"4A",x"66",x"DA",x"4A", -- 0x0A18
    x"66",x"DA",x"A6",x"DA",x"4C",x"2B",x"CA",x"E9", -- 0x0A20
    x"74",x"49",x"20",x"8C",x"00",x"FE",x"8D",x"01", -- 0x0A28
    x"FE",x"C8",x"8C",x"00",x"FE",x"8E",x"01",x"FE", -- 0x0A30
    x"60",x"20",x"81",x"CA",x"A2",x"1C",x"A0",x"2C", -- 0x0A38
    x"20",x"11",x"D4",x"0D",x"2D",x"03",x"30",x"39", -- 0x0A40
    x"A2",x"20",x"20",x"49",x"D1",x"A2",x"1C",x"20", -- 0x0A48
    x"49",x"D1",x"AD",x"1F",x"03",x"0D",x"1D",x"03", -- 0x0A50
    x"30",x"27",x"AD",x"23",x"03",x"D0",x"22",x"AE", -- 0x0A58
    x"55",x"03",x"AD",x"21",x"03",x"85",x"DA",x"AD", -- 0x0A60
    x"20",x"03",x"46",x"DA",x"6A",x"46",x"DA",x"D0", -- 0x0A68
    x"10",x"6A",x"4A",x"DD",x"EF",x"C3",x"F0",x"02", -- 0x0A70
    x"10",x"07",x"A0",x"00",x"A2",x"1C",x"20",x"7C", -- 0x0A78
    x"D4",x"A2",x"10",x"A0",x"28",x"4C",x"E6",x"CD", -- 0x0A80
    x"C8",x"98",x"A0",x"00",x"8C",x"4D",x"03",x"8D", -- 0x0A88
    x"4C",x"03",x"AD",x"4F",x"03",x"4A",x"F0",x"09", -- 0x0A90
    x"0E",x"4C",x"03",x"2E",x"4D",x"03",x"4A",x"90", -- 0x0A98
    x"F7",x"60",x"A2",x"20",x"A0",x"0C",x"20",x"8A", -- 0x0AA0
    x"D4",x"4C",x"B8",x"D1",x"20",x"C5",x"C5",x"20", -- 0x0AA8
    x"88",x"C5",x"D0",x"13",x"AE",x"60",x"03",x"F0", -- 0x0AB0
    x"09",x"85",x"DE",x"A9",x"C0",x"85",x"DF",x"4C", -- 0x0AB8
    x"BF",x"CF",x"A9",x"20",x"4C",x"DC",x"CF",x"A9", -- 0x0AC0
    x"7F",x"20",x"3E",x"D0",x"AE",x"5A",x"03",x"A0", -- 0x0AC8
    x"00",x"4C",x"63",x"CF",x"48",x"8A",x"18",x"6D", -- 0x0AD0
    x"52",x"03",x"AA",x"68",x"6D",x"53",x"03",x"60", -- 0x0AD8
    x"20",x"14",x"CB",x"20",x"D9",x"E9",x"90",x"02", -- 0x0AE0
    x"30",x"F6",x"A5",x"D0",x"49",x"04",x"29",x"46", -- 0x0AE8
    x"D0",x"2A",x"AD",x"69",x"02",x"30",x"22",x"AD", -- 0x0AF0
    x"19",x"03",x"CD",x"09",x"03",x"90",x"1A",x"4A", -- 0x0AF8
    x"4A",x"38",x"6D",x"69",x"02",x"6D",x"0B",x"03", -- 0x0B00
    x"CD",x"09",x"03",x"90",x"0C",x"18",x"20",x"D9", -- 0x0B08
    x"E9",x"38",x"10",x"FA",x"A9",x"FF",x"8D",x"69", -- 0x0B10
    x"02",x"EE",x"69",x"02",x"60",x"48",x"A2",x"7F", -- 0x0B18
    x"A9",x"00",x"85",x"D0",x"9D",x"FF",x"02",x"CA", -- 0x0B20
    x"D0",x"FA",x"20",x"07",x"CD",x"68",x"A2",x"7F", -- 0x0B28
    x"8E",x"66",x"03",x"2C",x"8E",x"02",x"30",x"02", -- 0x0B30
    x"09",x"04",x"29",x"07",x"AA",x"8E",x"55",x"03", -- 0x0B38
    x"BD",x"14",x"C4",x"8D",x"60",x"03",x"BD",x"FF", -- 0x0B40
    x"C3",x"8D",x"4F",x"03",x"BD",x"3A",x"C4",x"8D", -- 0x0B48
    x"61",x"03",x"D0",x"02",x"A9",x"07",x"0A",x"A8", -- 0x0B50
    x"B9",x"06",x"C4",x"8D",x"63",x"03",x"0A",x"10", -- 0x0B58
    x"FD",x"8D",x"62",x"03",x"BC",x"40",x"C4",x"8C", -- 0x0B60
    x"56",x"03",x"B9",x"4F",x"C4",x"20",x"F8",x"E9", -- 0x0B68
    x"B9",x"4B",x"C4",x"20",x"F8",x"E9",x"B9",x"59", -- 0x0B70
    x"C4",x"8D",x"54",x"03",x"B9",x"5E",x"C4",x"8D", -- 0x0B78
    x"4E",x"03",x"98",x"69",x"02",x"49",x"07",x"4A", -- 0x0B80
    x"AA",x"BD",x"66",x"C4",x"85",x"E0",x"A9",x"C3", -- 0x0B88
    x"85",x"E1",x"BD",x"63",x"C4",x"8D",x"52",x"03", -- 0x0B90
    x"8E",x"53",x"03",x"A9",x"43",x"20",x"A8",x"C5", -- 0x0B98
    x"AE",x"55",x"03",x"BD",x"F7",x"C3",x"20",x"00", -- 0x0BA0
    x"EA",x"08",x"78",x"BE",x"69",x"C4",x"A0",x"0B", -- 0x0BA8
    x"BD",x"6E",x"C4",x"20",x"5E",x"C9",x"CA",x"88", -- 0x0BB0
    x"10",x"F6",x"28",x"20",x"39",x"C8",x"20",x"BD", -- 0x0BB8
    x"C9",x"A2",x"00",x"AD",x"4E",x"03",x"8E",x"50", -- 0x0BC0
    x"03",x"8D",x"51",x"03",x"20",x"F6",x"C9",x"A0", -- 0x0BC8
    x"0C",x"20",x"2B",x"CA",x"AD",x"58",x"03",x"AE", -- 0x0BD0
    x"56",x"03",x"BC",x"54",x"C4",x"8C",x"5D",x"03", -- 0x0BD8
    x"A0",x"CC",x"8C",x"5E",x"03",x"A2",x"00",x"8E", -- 0x0BE0
    x"69",x"02",x"8E",x"18",x"03",x"8E",x"19",x"03", -- 0x0BE8
    x"6C",x"5D",x"03",x"20",x"3E",x"D0",x"A0",x"00", -- 0x0BF0
    x"B1",x"DE",x"C8",x"91",x"F0",x"C0",x"08",x"D0", -- 0x0BF8
    x"F7",x"60",x"9D",x"00",x"30",x"9D",x"00",x"31", -- 0x0C00
    x"9D",x"00",x"32",x"9D",x"00",x"33",x"9D",x"00", -- 0x0C08
    x"34",x"9D",x"00",x"35",x"9D",x"00",x"36",x"9D", -- 0x0C10
    x"00",x"37",x"9D",x"00",x"38",x"9D",x"00",x"39", -- 0x0C18
    x"9D",x"00",x"3A",x"9D",x"00",x"3B",x"9D",x"00", -- 0x0C20
    x"3C",x"9D",x"00",x"3D",x"9D",x"00",x"3E",x"9D", -- 0x0C28
    x"00",x"3F",x"9D",x"00",x"40",x"9D",x"00",x"41", -- 0x0C30
    x"9D",x"00",x"42",x"9D",x"00",x"43",x"9D",x"00", -- 0x0C38
    x"44",x"9D",x"00",x"45",x"9D",x"00",x"46",x"9D", -- 0x0C40
    x"00",x"47",x"9D",x"00",x"48",x"9D",x"00",x"49", -- 0x0C48
    x"9D",x"00",x"4A",x"9D",x"00",x"4B",x"9D",x"00", -- 0x0C50
    x"4C",x"9D",x"00",x"4D",x"9D",x"00",x"4E",x"9D", -- 0x0C58
    x"00",x"4F",x"9D",x"00",x"50",x"9D",x"00",x"51", -- 0x0C60
    x"9D",x"00",x"52",x"9D",x"00",x"53",x"9D",x"00", -- 0x0C68
    x"54",x"9D",x"00",x"55",x"9D",x"00",x"56",x"9D", -- 0x0C70
    x"00",x"57",x"9D",x"00",x"58",x"9D",x"00",x"59", -- 0x0C78
    x"9D",x"00",x"5A",x"9D",x"00",x"5B",x"9D",x"00", -- 0x0C80
    x"5C",x"9D",x"00",x"5D",x"9D",x"00",x"5E",x"9D", -- 0x0C88
    x"00",x"5F",x"9D",x"00",x"60",x"9D",x"00",x"61", -- 0x0C90
    x"9D",x"00",x"62",x"9D",x"00",x"63",x"9D",x"00", -- 0x0C98
    x"64",x"9D",x"00",x"65",x"9D",x"00",x"66",x"9D", -- 0x0CA0
    x"00",x"67",x"9D",x"00",x"68",x"9D",x"00",x"69", -- 0x0CA8
    x"9D",x"00",x"6A",x"9D",x"00",x"6B",x"9D",x"00", -- 0x0CB0
    x"6C",x"9D",x"00",x"6D",x"9D",x"00",x"6E",x"9D", -- 0x0CB8
    x"00",x"6F",x"9D",x"00",x"70",x"9D",x"00",x"71", -- 0x0CC0
    x"9D",x"00",x"72",x"9D",x"00",x"73",x"9D",x"00", -- 0x0CC8
    x"74",x"9D",x"00",x"75",x"9D",x"00",x"76",x"9D", -- 0x0CD0
    x"00",x"77",x"9D",x"00",x"78",x"9D",x"00",x"79", -- 0x0CD8
    x"9D",x"00",x"7A",x"9D",x"00",x"7B",x"9D",x"00", -- 0x0CE0
    x"7C",x"9D",x"00",x"7D",x"9D",x"00",x"7E",x"9D", -- 0x0CE8
    x"00",x"7F",x"E8",x"F0",x"70",x"6C",x"5D",x"03", -- 0x0CF0
    x"48",x"8A",x"38",x"ED",x"52",x"03",x"AA",x"68", -- 0x0CF8
    x"ED",x"53",x"03",x"CD",x"4E",x"03",x"60",x"A9", -- 0x0D00
    x"0F",x"8D",x"67",x"03",x"A9",x"0C",x"A0",x"06", -- 0x0D08
    x"99",x"68",x"03",x"88",x"10",x"FA",x"E0",x"07", -- 0x0D10
    x"90",x"02",x"A2",x"06",x"8E",x"46",x"02",x"AD", -- 0x0D18
    x"43",x"02",x"A2",x"00",x"EC",x"46",x"02",x"B0", -- 0x0D20
    x"0B",x"BC",x"BA",x"C4",x"99",x"68",x"03",x"69", -- 0x0D28
    x"01",x"E8",x"D0",x"F0",x"8D",x"44",x"02",x"A8", -- 0x0D30
    x"F0",x"CC",x"A2",x"11",x"4C",x"68",x"F1",x"A9", -- 0x0D38
    x"02",x"24",x"D0",x"D0",x"02",x"50",x"32",x"AD", -- 0x0D40
    x"09",x"03",x"90",x"03",x"AD",x"0B",x"03",x"70", -- 0x0D48
    x"08",x"8D",x"19",x"03",x"68",x"68",x"4C",x"AF", -- 0x0D50
    x"C6",x"08",x"CD",x"65",x"03",x"F0",x"19",x"28", -- 0x0D58
    x"90",x"04",x"CE",x"65",x"03",x"60",x"EE",x"65", -- 0x0D60
    x"03",x"60",x"08",x"48",x"AC",x"4F",x"03",x"88", -- 0x0D68
    x"D0",x"1D",x"AD",x"38",x"03",x"91",x"D8",x"68", -- 0x0D70
    x"28",x"60",x"08",x"48",x"AC",x"4F",x"03",x"88", -- 0x0D78
    x"D0",x"0D",x"B1",x"D8",x"8D",x"38",x"03",x"AD", -- 0x0D80
    x"66",x"03",x"91",x"D8",x"4C",x"77",x"CD",x"A9", -- 0x0D88
    x"FF",x"C0",x"1F",x"D0",x"02",x"A9",x"3F",x"85", -- 0x0D90
    x"DA",x"B1",x"D8",x"45",x"DA",x"91",x"D8",x"88", -- 0x0D98
    x"10",x"F7",x"30",x"D3",x"20",x"5B",x"CE",x"AD", -- 0x0DA0
    x"09",x"03",x"8D",x"19",x"03",x"20",x"06",x"CF", -- 0x0DA8
    x"20",x"F8",x"CC",x"B0",x"03",x"6D",x"54",x"03", -- 0x0DB0
    x"85",x"DB",x"86",x"DA",x"85",x"DC",x"B0",x"06", -- 0x0DB8
    x"20",x"73",x"CE",x"4C",x"CE",x"CD",x"20",x"F8", -- 0x0DC0
    x"CC",x"90",x"F5",x"20",x"38",x"CE",x"A5",x"DC", -- 0x0DC8
    x"A6",x"DA",x"85",x"D9",x"86",x"D8",x"C6",x"DE", -- 0x0DD0
    x"D0",x"D6",x"A2",x"28",x"A0",x"18",x"A9",x"02", -- 0x0DD8
    x"D0",x"06",x"A2",x"24",x"A0",x"14",x"A9",x"04", -- 0x0DE0
    x"85",x"DA",x"BD",x"00",x"03",x"48",x"B9",x"00", -- 0x0DE8
    x"03",x"9D",x"00",x"03",x"68",x"99",x"00",x"03", -- 0x0DF0
    x"E8",x"C8",x"C6",x"DA",x"D0",x"EC",x"60",x"20", -- 0x0DF8
    x"5B",x"CE",x"AC",x"0B",x"03",x"8C",x"19",x"03", -- 0x0E00
    x"20",x"06",x"CF",x"20",x"D4",x"CA",x"10",x"04", -- 0x0E08
    x"38",x"ED",x"54",x"03",x"85",x"DB",x"86",x"DA", -- 0x0E10
    x"85",x"DC",x"90",x"06",x"20",x"73",x"CE",x"4C", -- 0x0E18
    x"2A",x"CE",x"20",x"D4",x"CA",x"30",x"F5",x"20", -- 0x0E20
    x"38",x"CE",x"A5",x"DC",x"A6",x"DA",x"85",x"D9", -- 0x0E28
    x"86",x"D8",x"C6",x"DE",x"D0",x"D5",x"F0",x"A2", -- 0x0E30
    x"AE",x"4D",x"03",x"F0",x"10",x"A0",x"00",x"B1", -- 0x0E38
    x"DA",x"91",x"D8",x"C8",x"D0",x"F9",x"E6",x"D9", -- 0x0E40
    x"E6",x"DB",x"CA",x"D0",x"F2",x"AC",x"4C",x"03", -- 0x0E48
    x"F0",x"08",x"88",x"B1",x"DA",x"91",x"D8",x"98", -- 0x0E50
    x"D0",x"F8",x"60",x"20",x"DA",x"CD",x"38",x"AD", -- 0x0E58
    x"09",x"03",x"ED",x"0B",x"03",x"85",x"DE",x"D0", -- 0x0E60
    x"05",x"68",x"68",x"4C",x"DA",x"CD",x"AD",x"08", -- 0x0E68
    x"03",x"10",x"70",x"A5",x"DA",x"48",x"38",x"AD", -- 0x0E70
    x"0A",x"03",x"ED",x"08",x"03",x"85",x"DF",x"AC", -- 0x0E78
    x"4F",x"03",x"88",x"B1",x"DA",x"91",x"D8",x"88", -- 0x0E80
    x"10",x"F9",x"A2",x"02",x"18",x"B5",x"D8",x"6D", -- 0x0E88
    x"4F",x"03",x"95",x"D8",x"B5",x"D9",x"69",x"00", -- 0x0E90
    x"10",x"04",x"38",x"ED",x"54",x"03",x"95",x"D9", -- 0x0E98
    x"CA",x"CA",x"F0",x"E8",x"C6",x"DF",x"10",x"D7", -- 0x0EA0
    x"68",x"85",x"DA",x"60",x"AD",x"18",x"03",x"48", -- 0x0EA8
    x"20",x"6E",x"CE",x"20",x"06",x"CF",x"38",x"AD", -- 0x0EB0
    x"0A",x"03",x"ED",x"08",x"03",x"85",x"DC",x"AD", -- 0x0EB8
    x"58",x"03",x"AC",x"4F",x"03",x"88",x"91",x"D8", -- 0x0EC0
    x"D0",x"FB",x"8A",x"18",x"6D",x"4F",x"03",x"AA", -- 0x0EC8
    x"A5",x"D9",x"69",x"00",x"10",x"04",x"38",x"ED", -- 0x0ED0
    x"54",x"03",x"86",x"D8",x"85",x"D9",x"C6",x"DC", -- 0x0ED8
    x"10",x"DD",x"68",x"8D",x"18",x"03",x"38",x"60", -- 0x0EE0
    x"AE",x"18",x"03",x"EC",x"08",x"03",x"30",x"F6", -- 0x0EE8
    x"EC",x"0A",x"03",x"F0",x"02",x"10",x"EF",x"AE", -- 0x0EF0
    x"19",x"03",x"EC",x"0B",x"03",x"30",x"E7",x"EC", -- 0x0EF8
    x"09",x"03",x"F0",x"02",x"10",x"E0",x"AD",x"19", -- 0x0F00
    x"03",x"0A",x"A8",x"B1",x"E0",x"85",x"D9",x"C8", -- 0x0F08
    x"A9",x"02",x"2D",x"56",x"03",x"08",x"B1",x"E0", -- 0x0F10
    x"28",x"F0",x"03",x"46",x"D9",x"6A",x"6D",x"50", -- 0x0F18
    x"03",x"85",x"D8",x"A5",x"D9",x"6D",x"51",x"03", -- 0x0F20
    x"A8",x"AD",x"18",x"03",x"AE",x"4F",x"03",x"CA", -- 0x0F28
    x"F0",x"12",x"E0",x"0F",x"F0",x"03",x"90",x"02", -- 0x0F30
    x"0A",x"0A",x"0A",x"0A",x"90",x"02",x"C8",x"C8", -- 0x0F38
    x"0A",x"90",x"02",x"C8",x"18",x"65",x"D8",x"85", -- 0x0F40
    x"D8",x"8D",x"4A",x"03",x"AA",x"98",x"69",x"00", -- 0x0F48
    x"8D",x"4B",x"03",x"10",x"04",x"38",x"ED",x"54", -- 0x0F50
    x"03",x"85",x"D9",x"18",x"60",x"AE",x"59",x"03", -- 0x0F58
    x"AC",x"5B",x"03",x"20",x"B3",x"D0",x"20",x"86", -- 0x0F60
    x"D4",x"A0",x"00",x"84",x"DC",x"A4",x"DC",x"B1", -- 0x0F68
    x"DE",x"F0",x"13",x"85",x"DD",x"10",x"03",x"20", -- 0x0F70
    x"E3",x"D0",x"EE",x"24",x"03",x"D0",x"03",x"EE", -- 0x0F78
    x"25",x"03",x"06",x"DD",x"D0",x"EF",x"A2",x"28", -- 0x0F80
    x"A0",x"24",x"20",x"82",x"D4",x"AC",x"26",x"03", -- 0x0F88
    x"D0",x"03",x"CE",x"27",x"03",x"CE",x"26",x"03", -- 0x0F90
    x"A4",x"DC",x"C8",x"C0",x"08",x"D0",x"CC",x"A2", -- 0x0F98
    x"28",x"A0",x"24",x"4C",x"8A",x"D4",x"A2",x"06", -- 0x0FA0
    x"A0",x"26",x"20",x"82",x"D4",x"A2",x"00",x"A0", -- 0x0FA8
    x"24",x"20",x"82",x"D4",x"4C",x"B8",x"D1",x"AE", -- 0x0FB0
    x"60",x"03",x"F0",x"20",x"20",x"3E",x"D0",x"AE", -- 0x0FB8
    x"60",x"03",x"A5",x"D0",x"29",x"20",x"D0",x"95", -- 0x0FC0
    x"A0",x"07",x"E0",x"03",x"F0",x"20",x"B0",x"4E", -- 0x0FC8
    x"B1",x"DE",x"05",x"D2",x"45",x"D3",x"91",x"D8", -- 0x0FD0
    x"88",x"10",x"F5",x"60",x"A0",x"02",x"D9",x"B6", -- 0x0FD8
    x"C4",x"F0",x"06",x"88",x"10",x"F8",x"81",x"D8", -- 0x0FE0
    x"60",x"B9",x"B7",x"C4",x"D0",x"F8",x"B1",x"DE", -- 0x0FE8
    x"48",x"4A",x"4A",x"4A",x"4A",x"AA",x"BD",x"1F", -- 0x0FF0
    x"C3",x"05",x"D2",x"45",x"D3",x"91",x"D8",x"98", -- 0x0FF8
    x"18",x"69",x"08",x"A8",x"68",x"29",x"0F",x"AA", -- 0x1000
    x"BD",x"1F",x"C3",x"05",x"D2",x"45",x"D3",x"91", -- 0x1008
    x"D8",x"98",x"E9",x"08",x"A8",x"10",x"D7",x"60", -- 0x1010
    x"98",x"E9",x"21",x"30",x"FA",x"A8",x"B1",x"DE", -- 0x1018
    x"85",x"DC",x"38",x"A9",x"00",x"26",x"DC",x"F0", -- 0x1020
    x"EF",x"2A",x"06",x"DC",x"2A",x"AA",x"BD",x"2F", -- 0x1028
    x"C3",x"05",x"D2",x"45",x"D3",x"91",x"D8",x"18", -- 0x1030
    x"98",x"69",x"08",x"A8",x"90",x"E5",x"0A",x"2A", -- 0x1038
    x"2A",x"85",x"DE",x"29",x"03",x"2A",x"AA",x"29", -- 0x1040
    x"03",x"69",x"BF",x"A8",x"BD",x"0D",x"C4",x"2C", -- 0x1048
    x"67",x"03",x"F0",x"03",x"BC",x"67",x"03",x"84", -- 0x1050
    x"DF",x"A5",x"DE",x"29",x"F8",x"85",x"DE",x"60", -- 0x1058
    x"A2",x"20",x"20",x"4D",x"D1",x"AD",x"1F",x"03", -- 0x1060
    x"C9",x"04",x"F0",x"6D",x"A0",x"05",x"29",x"03", -- 0x1068
    x"F0",x"0E",x"4A",x"B0",x"03",x"88",x"D0",x"08", -- 0x1070
    x"AA",x"BC",x"5B",x"03",x"BD",x"59",x"03",x"AA", -- 0x1078
    x"20",x"B3",x"D0",x"AD",x"1F",x"03",x"30",x"23", -- 0x1080
    x"0A",x"10",x"3B",x"29",x"F0",x"0A",x"F0",x"46", -- 0x1088
    x"49",x"40",x"F0",x"14",x"48",x"20",x"DC",x"D0", -- 0x1090
    x"68",x"49",x"60",x"F0",x"11",x"C9",x"40",x"D0", -- 0x1098
    x"0A",x"A9",x"02",x"85",x"DC",x"4C",x"06",x"D5", -- 0x10A0
    x"4C",x"EA",x"D5",x"4C",x"38",x"C9",x"85",x"DC", -- 0x10A8
    x"4C",x"BF",x"D4",x"8A",x"19",x"1C",x"C4",x"59", -- 0x10B0
    x"1D",x"C4",x"85",x"D4",x"8A",x"19",x"1B",x"C4", -- 0x10B8
    x"59",x"20",x"C4",x"85",x"D5",x"60",x"0A",x"30", -- 0x10C0
    x"E2",x"0A",x"0A",x"10",x"03",x"20",x"EB",x"D0", -- 0x10C8
    x"20",x"ED",x"D1",x"4C",x"D9",x"D0",x"20",x"EB", -- 0x10D0
    x"D0",x"20",x"E2",x"CD",x"A0",x"24",x"A2",x"20", -- 0x10D8
    x"4C",x"8A",x"D4",x"A2",x"24",x"20",x"5F",x"D8", -- 0x10E0
    x"F0",x"06",x"60",x"20",x"5D",x"D8",x"D0",x"13", -- 0x10E8
    x"AC",x"1A",x"03",x"A5",x"D1",x"25",x"D4",x"11", -- 0x10F0
    x"D6",x"85",x"DA",x"A5",x"D5",x"25",x"D1",x"45", -- 0x10F8
    x"DA",x"91",x"D6",x"60",x"B1",x"D6",x"05",x"D4", -- 0x1100
    x"45",x"D5",x"91",x"D6",x"60",x"A2",x"24",x"A0", -- 0x1108
    x"00",x"84",x"DA",x"A0",x"02",x"20",x"28",x"D1", -- 0x1110
    x"06",x"DA",x"06",x"DA",x"CA",x"CA",x"A0",x"00", -- 0x1118
    x"20",x"28",x"D1",x"E8",x"E8",x"A5",x"DA",x"60", -- 0x1120
    x"BD",x"02",x"03",x"D9",x"00",x"03",x"BD",x"03", -- 0x1128
    x"03",x"F9",x"01",x"03",x"30",x"10",x"B9",x"04", -- 0x1130
    x"03",x"DD",x"02",x"03",x"B9",x"05",x"03",x"FD", -- 0x1138
    x"03",x"03",x"10",x"04",x"E6",x"DA",x"E6",x"DA", -- 0x1140
    x"60",x"A9",x"FF",x"D0",x"03",x"AD",x"1F",x"03", -- 0x1148
    x"85",x"DA",x"A0",x"02",x"20",x"76",x"D1",x"20", -- 0x1150
    x"AD",x"D1",x"A0",x"00",x"CA",x"CA",x"20",x"76", -- 0x1158
    x"D1",x"AC",x"61",x"03",x"C0",x"03",x"F0",x"05", -- 0x1160
    x"B0",x"06",x"20",x"AD",x"D1",x"20",x"AD",x"D1", -- 0x1168
    x"AD",x"56",x"03",x"D0",x"38",x"60",x"18",x"A5", -- 0x1170
    x"DA",x"29",x"04",x"F0",x"09",x"BD",x"02",x"03", -- 0x1178
    x"48",x"BD",x"03",x"03",x"90",x"0E",x"BD",x"02", -- 0x1180
    x"03",x"79",x"10",x"03",x"48",x"BD",x"03",x"03", -- 0x1188
    x"79",x"11",x"03",x"18",x"99",x"11",x"03",x"79", -- 0x1190
    x"0D",x"03",x"9D",x"03",x"03",x"68",x"99",x"10", -- 0x1198
    x"03",x"18",x"79",x"0C",x"03",x"9D",x"02",x"03", -- 0x11A0
    x"90",x"03",x"FE",x"03",x"03",x"BD",x"03",x"03", -- 0x11A8
    x"0A",x"7E",x"03",x"03",x"7E",x"02",x"03",x"60", -- 0x11B0
    x"A0",x"10",x"20",x"88",x"D4",x"A2",x"02",x"A0", -- 0x11B8
    x"02",x"20",x"D5",x"D1",x"A2",x"00",x"A0",x"04", -- 0x11C0
    x"AD",x"61",x"03",x"88",x"4A",x"D0",x"FC",x"AD", -- 0x11C8
    x"56",x"03",x"F0",x"01",x"C8",x"1E",x"10",x"03", -- 0x11D0
    x"3E",x"11",x"03",x"88",x"D0",x"F7",x"38",x"20", -- 0x11D8
    x"E3",x"D1",x"E8",x"BD",x"10",x"03",x"FD",x"0C", -- 0x11E0
    x"03",x"9D",x"10",x"03",x"60",x"20",x"0D",x"D4", -- 0x11E8
    x"AD",x"2B",x"03",x"4D",x"29",x"03",x"30",x"0F", -- 0x11F0
    x"AD",x"2A",x"03",x"CD",x"28",x"03",x"AD",x"2B", -- 0x11F8
    x"03",x"ED",x"29",x"03",x"4C",x"14",x"D2",x"AD", -- 0x1200
    x"28",x"03",x"18",x"6D",x"2A",x"03",x"AD",x"29", -- 0x1208
    x"03",x"6D",x"2B",x"03",x"6A",x"A2",x"00",x"4D", -- 0x1210
    x"2B",x"03",x"10",x"02",x"A2",x"02",x"86",x"DE", -- 0x1218
    x"BD",x"AA",x"C4",x"8D",x"5D",x"03",x"BD",x"AB", -- 0x1220
    x"C4",x"8D",x"5E",x"03",x"BD",x"29",x"03",x"10", -- 0x1228
    x"04",x"A2",x"24",x"D0",x"02",x"A2",x"20",x"86", -- 0x1230
    x"DF",x"A0",x"2C",x"20",x"8A",x"D4",x"A5",x"DF", -- 0x1238
    x"49",x"04",x"85",x"DD",x"05",x"DE",x"AA",x"20", -- 0x1240
    x"80",x"D4",x"AD",x"1F",x"03",x"29",x"10",x"0A", -- 0x1248
    x"0A",x"0A",x"85",x"DB",x"A2",x"2C",x"20",x"0F", -- 0x1250
    x"D1",x"85",x"DC",x"F0",x"06",x"A9",x"40",x"05", -- 0x1258
    x"DB",x"85",x"DB",x"A6",x"DD",x"20",x"0F",x"D1", -- 0x1260
    x"24",x"DC",x"F0",x"01",x"60",x"A6",x"DE",x"F0", -- 0x1268
    x"02",x"4A",x"4A",x"29",x"02",x"F0",x"07",x"8A", -- 0x1270
    x"09",x"04",x"AA",x"20",x"80",x"D4",x"20",x"2C", -- 0x1278
    x"D4",x"A5",x"DE",x"49",x"02",x"AA",x"A8",x"AD", -- 0x1280
    x"29",x"03",x"4D",x"2B",x"03",x"10",x"01",x"E8", -- 0x1288
    x"BD",x"AE",x"C4",x"8D",x"32",x"03",x"BD",x"B2", -- 0x1290
    x"C4",x"8D",x"33",x"03",x"A9",x"7F",x"8D",x"34", -- 0x1298
    x"03",x"24",x"DB",x"70",x"29",x"BD",x"47",x"C4", -- 0x12A0
    x"AA",x"38",x"BD",x"00",x"03",x"F9",x"2C",x"03", -- 0x12A8
    x"85",x"DA",x"BD",x"01",x"03",x"F9",x"2D",x"03", -- 0x12B0
    x"A4",x"DA",x"AA",x"10",x"03",x"20",x"9B",x"D4", -- 0x12B8
    x"AA",x"C8",x"D0",x"01",x"E8",x"8A",x"F0",x"02", -- 0x12C0
    x"A0",x"00",x"84",x"DF",x"F0",x"09",x"8A",x"4A", -- 0x12C8
    x"6A",x"09",x"02",x"45",x"DE",x"85",x"DE",x"A2", -- 0x12D0
    x"2C",x"20",x"64",x"D8",x"A6",x"DC",x"D0",x"02", -- 0x12D8
    x"C6",x"DD",x"CA",x"A5",x"DB",x"F0",x"1F",x"10", -- 0x12E0
    x"10",x"2C",x"34",x"03",x"10",x"05",x"CE",x"34", -- 0x12E8
    x"03",x"D0",x"23",x"EE",x"34",x"03",x"0A",x"10", -- 0x12F0
    x"0D",x"86",x"DC",x"A2",x"2C",x"20",x"5F",x"D8", -- 0x12F8
    x"A6",x"DC",x"09",x"00",x"D0",x"10",x"A5",x"D1", -- 0x1300
    x"25",x"D4",x"11",x"D6",x"85",x"DA",x"A5",x"D5", -- 0x1308
    x"25",x"D1",x"45",x"DA",x"91",x"D6",x"38",x"AD", -- 0x1310
    x"35",x"03",x"ED",x"37",x"03",x"8D",x"35",x"03", -- 0x1318
    x"AD",x"36",x"03",x"ED",x"38",x"03",x"B0",x"11", -- 0x1320
    x"85",x"DA",x"AD",x"35",x"03",x"6D",x"39",x"03", -- 0x1328
    x"8D",x"35",x"03",x"A5",x"DA",x"6D",x"3A",x"03", -- 0x1330
    x"18",x"8D",x"36",x"03",x"08",x"B0",x"09",x"6C", -- 0x1338
    x"32",x"03",x"88",x"10",x"03",x"20",x"D3",x"D3", -- 0x1340
    x"6C",x"5D",x"03",x"C8",x"C0",x"08",x"D0",x"F8", -- 0x1348
    x"18",x"A5",x"D6",x"6D",x"52",x"03",x"85",x"D6", -- 0x1350
    x"A5",x"D7",x"6D",x"53",x"03",x"10",x"04",x"38", -- 0x1358
    x"ED",x"54",x"03",x"85",x"D7",x"A0",x"00",x"6C", -- 0x1360
    x"5D",x"03",x"46",x"D1",x"90",x"DA",x"20",x"ED", -- 0x1368
    x"D3",x"6C",x"5D",x"03",x"06",x"D1",x"90",x"D0", -- 0x1370
    x"20",x"FD",x"D3",x"6C",x"5D",x"03",x"88",x"10", -- 0x1378
    x"0C",x"20",x"D3",x"D3",x"D0",x"07",x"46",x"D1", -- 0x1380
    x"90",x"03",x"20",x"ED",x"D3",x"28",x"E8",x"D0", -- 0x1388
    x"04",x"E6",x"DD",x"F0",x"0A",x"24",x"DB",x"70", -- 0x1390
    x"07",x"B0",x"35",x"C6",x"DF",x"D0",x"31",x"60", -- 0x1398
    x"A5",x"DE",x"86",x"DC",x"29",x"02",x"AA",x"B0", -- 0x13A0
    x"19",x"24",x"DE",x"30",x"0A",x"FE",x"2C",x"03", -- 0x13A8
    x"D0",x"10",x"FE",x"2D",x"03",x"90",x"0B",x"BD", -- 0x13B0
    x"2C",x"03",x"D0",x"03",x"DE",x"2D",x"03",x"DE", -- 0x13B8
    x"2C",x"03",x"8A",x"49",x"02",x"AA",x"FE",x"2C", -- 0x13C0
    x"03",x"D0",x"03",x"FE",x"2D",x"03",x"A6",x"DC", -- 0x13C8
    x"4C",x"E3",x"D2",x"38",x"A5",x"D6",x"ED",x"52", -- 0x13D0
    x"03",x"85",x"D6",x"A5",x"D7",x"ED",x"53",x"03", -- 0x13D8
    x"CD",x"4E",x"03",x"B0",x"03",x"6D",x"54",x"03", -- 0x13E0
    x"85",x"D7",x"A0",x"07",x"60",x"AD",x"62",x"03", -- 0x13E8
    x"85",x"D1",x"A5",x"D6",x"69",x"07",x"85",x"D6", -- 0x13F0
    x"90",x"02",x"E6",x"D7",x"60",x"AD",x"63",x"03", -- 0x13F8
    x"85",x"D1",x"A5",x"D6",x"D0",x"02",x"C6",x"D7", -- 0x1400
    x"E9",x"08",x"85",x"D6",x"60",x"A0",x"28",x"A2", -- 0x1408
    x"20",x"20",x"18",x"D4",x"E8",x"E8",x"C8",x"C8", -- 0x1410
    x"38",x"BD",x"04",x"03",x"FD",x"00",x"03",x"99", -- 0x1418
    x"00",x"03",x"BD",x"05",x"03",x"FD",x"01",x"03", -- 0x1420
    x"99",x"01",x"03",x"60",x"A5",x"DE",x"D0",x"07", -- 0x1428
    x"A2",x"28",x"A0",x"2A",x"20",x"DE",x"CD",x"A2", -- 0x1430
    x"28",x"A0",x"37",x"20",x"8A",x"D4",x"38",x"A6", -- 0x1438
    x"DE",x"AD",x"30",x"03",x"FD",x"2C",x"03",x"A8", -- 0x1440
    x"AD",x"31",x"03",x"FD",x"2D",x"03",x"30",x"03", -- 0x1448
    x"20",x"9B",x"D4",x"85",x"DD",x"84",x"DC",x"A2", -- 0x1450
    x"35",x"20",x"67",x"D4",x"4A",x"9D",x"01",x"03", -- 0x1458
    x"98",x"6A",x"9D",x"00",x"03",x"CA",x"CA",x"BC", -- 0x1460
    x"04",x"03",x"BD",x"05",x"03",x"10",x"0C",x"20", -- 0x1468
    x"9B",x"D4",x"9D",x"05",x"03",x"48",x"98",x"9D", -- 0x1470
    x"04",x"03",x"68",x"60",x"A9",x"08",x"D0",x"0C", -- 0x1478
    x"A0",x"30",x"A9",x"02",x"D0",x"06",x"A0",x"28", -- 0x1480
    x"A2",x"24",x"A9",x"04",x"85",x"DA",x"BD",x"00", -- 0x1488
    x"03",x"99",x"00",x"03",x"E8",x"C8",x"C6",x"DA", -- 0x1490
    x"D0",x"F4",x"60",x"48",x"98",x"49",x"FF",x"A8", -- 0x1498
    x"68",x"49",x"FF",x"C8",x"D0",x"03",x"18",x"69", -- 0x14A0
    x"01",x"60",x"20",x"5D",x"D8",x"D0",x"08",x"B1", -- 0x14A8
    x"D6",x"4D",x"5A",x"03",x"85",x"DA",x"60",x"68", -- 0x14B0
    x"68",x"EE",x"26",x"03",x"4C",x"45",x"D5",x"20", -- 0x14B8
    x"AA",x"D4",x"25",x"D1",x"D0",x"F3",x"A2",x"00", -- 0x14C0
    x"20",x"92",x"D5",x"F0",x"2D",x"AC",x"1A",x"03", -- 0x14C8
    x"06",x"D1",x"B0",x"05",x"20",x"74",x"D5",x"90", -- 0x14D0
    x"21",x"20",x"FD",x"D3",x"B1",x"D6",x"4D",x"5A", -- 0x14D8
    x"03",x"85",x"DA",x"D0",x"12",x"38",x"8A",x"6D", -- 0x14E0
    x"61",x"03",x"90",x"04",x"E6",x"DB",x"10",x"07", -- 0x14E8
    x"AA",x"20",x"04",x"D1",x"38",x"B0",x"E2",x"20", -- 0x14F0
    x"74",x"D5",x"A0",x"00",x"20",x"AC",x"D5",x"A0", -- 0x14F8
    x"20",x"A2",x"24",x"20",x"E6",x"CD",x"20",x"AA", -- 0x1500
    x"D4",x"A2",x"04",x"20",x"92",x"D5",x"8A",x"D0", -- 0x1508
    x"02",x"C6",x"DB",x"CA",x"20",x"4B",x"D5",x"90", -- 0x1510
    x"27",x"20",x"ED",x"D3",x"B1",x"D6",x"4D",x"5A", -- 0x1518
    x"03",x"85",x"DA",x"A5",x"DC",x"D0",x"ED",x"A5", -- 0x1520
    x"DA",x"D0",x"12",x"38",x"8A",x"6D",x"61",x"03", -- 0x1528
    x"90",x"04",x"E6",x"DB",x"10",x"07",x"AA",x"20", -- 0x1530
    x"04",x"D1",x"38",x"B0",x"DC",x"20",x"4B",x"D5", -- 0x1538
    x"A0",x"04",x"20",x"AC",x"D5",x"20",x"D9",x"D0", -- 0x1540
    x"4C",x"B8",x"D1",x"A5",x"D1",x"48",x"18",x"90", -- 0x1548
    x"0F",x"68",x"E8",x"D0",x"04",x"E6",x"DB",x"10", -- 0x1550
    x"16",x"46",x"D1",x"B0",x"12",x"05",x"D1",x"48", -- 0x1558
    x"A5",x"D1",x"24",x"DA",x"08",x"68",x"45",x"DC", -- 0x1560
    x"48",x"28",x"F0",x"E5",x"68",x"45",x"D1",x"85", -- 0x1568
    x"D1",x"4C",x"F0",x"D0",x"A9",x"00",x"18",x"90", -- 0x1570
    x"0A",x"E8",x"D0",x"04",x"E6",x"DB",x"10",x"EF", -- 0x1578
    x"0A",x"B0",x"0B",x"05",x"D1",x"24",x"DA",x"F0", -- 0x1580
    x"F0",x"45",x"D1",x"4A",x"90",x"E1",x"6A",x"38", -- 0x1588
    x"B0",x"DD",x"BD",x"00",x"03",x"38",x"ED",x"20", -- 0x1590
    x"03",x"A8",x"BD",x"01",x"03",x"ED",x"21",x"03", -- 0x1598
    x"30",x"03",x"20",x"9B",x"D4",x"85",x"DB",x"98", -- 0x15A0
    x"AA",x"05",x"DB",x"60",x"84",x"DA",x"8A",x"A8", -- 0x15A8
    x"A5",x"DB",x"30",x"02",x"A9",x"00",x"A6",x"DA", -- 0x15B0
    x"D0",x"03",x"20",x"9B",x"D4",x"48",x"18",x"98", -- 0x15B8
    x"7D",x"00",x"03",x"8D",x"20",x"03",x"68",x"7D", -- 0x15C0
    x"01",x"03",x"8D",x"21",x"03",x"60",x"A9",x"03", -- 0x15C8
    x"20",x"D5",x"D5",x"A9",x"07",x"48",x"20",x"E2", -- 0x15D0
    x"CD",x"20",x"B8",x"D1",x"A2",x"03",x"68",x"A8", -- 0x15D8
    x"BD",x"10",x"03",x"91",x"F0",x"88",x"CA",x"10", -- 0x15E0
    x"F7",x"60",x"A2",x"20",x"A0",x"3E",x"20",x"7C", -- 0x15E8
    x"D4",x"20",x"32",x"D6",x"A2",x"14",x"A0",x"24", -- 0x15F0
    x"20",x"36",x"D6",x"20",x"32",x"D6",x"A2",x"20", -- 0x15F8
    x"A0",x"2A",x"20",x"11",x"D4",x"AD",x"2B",x"03", -- 0x1600
    x"8D",x"32",x"03",x"A2",x"28",x"20",x"59",x"D4", -- 0x1608
    x"A0",x"2E",x"20",x"DE",x"D0",x"20",x"E2",x"CD", -- 0x1610
    x"18",x"20",x"58",x"D6",x"20",x"E2",x"CD",x"A2", -- 0x1618
    x"20",x"20",x"E4",x"CD",x"38",x"20",x"58",x"D6", -- 0x1620
    x"A2",x"3E",x"A0",x"20",x"20",x"7C",x"D4",x"4C", -- 0x1628
    x"D9",x"D0",x"A2",x"20",x"A0",x"14",x"BD",x"02", -- 0x1630
    x"03",x"D9",x"02",x"03",x"BD",x"03",x"03",x"F9", -- 0x1638
    x"03",x"03",x"30",x"13",x"4C",x"E6",x"CD",x"AD", -- 0x1640
    x"18",x"03",x"38",x"ED",x"08",x"03",x"AA",x"AD", -- 0x1648
    x"19",x"03",x"38",x"ED",x"0B",x"03",x"A8",x"60", -- 0x1650
    x"08",x"A2",x"20",x"A0",x"35",x"20",x"11",x"D4", -- 0x1658
    x"AD",x"36",x"03",x"8D",x"3D",x"03",x"A2",x"33", -- 0x1660
    x"20",x"59",x"D4",x"A0",x"39",x"20",x"DE",x"D0", -- 0x1668
    x"38",x"AD",x"22",x"03",x"ED",x"26",x"03",x"8D", -- 0x1670
    x"1B",x"03",x"AD",x"23",x"03",x"ED",x"27",x"03", -- 0x1678
    x"8D",x"1C",x"03",x"0D",x"1B",x"03",x"F0",x"17", -- 0x1680
    x"20",x"A2",x"D6",x"A2",x"33",x"20",x"74",x"D7", -- 0x1688
    x"A2",x"28",x"20",x"74",x"D7",x"EE",x"1B",x"03", -- 0x1690
    x"D0",x"EE",x"EE",x"1C",x"03",x"D0",x"E9",x"28", -- 0x1698
    x"90",x"B5",x"A2",x"39",x"A0",x"2E",x"86",x"DE", -- 0x16A0
    x"BD",x"00",x"03",x"D9",x"00",x"03",x"BD",x"01", -- 0x16A8
    x"03",x"F9",x"01",x"03",x"30",x"06",x"98",x"A4", -- 0x16B0
    x"DE",x"AA",x"86",x"DE",x"84",x"DF",x"B9",x"00", -- 0x16B8
    x"03",x"48",x"B9",x"01",x"03",x"48",x"A6",x"DF", -- 0x16C0
    x"20",x"0F",x"D1",x"F0",x"0D",x"C9",x"02",x"D0", -- 0x16C8
    x"3D",x"A2",x"04",x"A4",x"DF",x"20",x"82",x"D4", -- 0x16D0
    x"A6",x"DF",x"20",x"64",x"D8",x"A6",x"DE",x"20", -- 0x16D8
    x"0F",x"D1",x"4A",x"D0",x"29",x"90",x"02",x"A2", -- 0x16E0
    x"00",x"A4",x"DF",x"38",x"B9",x"00",x"03",x"FD", -- 0x16E8
    x"00",x"03",x"85",x"DC",x"B9",x"01",x"03",x"FD", -- 0x16F0
    x"01",x"03",x"85",x"DD",x"A9",x"00",x"0A",x"05", -- 0x16F8
    x"D1",x"A4",x"DC",x"D0",x"14",x"C6",x"DD",x"10", -- 0x1700
    x"10",x"85",x"D1",x"20",x"F0",x"D0",x"A6",x"DF", -- 0x1708
    x"68",x"9D",x"01",x"03",x"68",x"9D",x"00",x"03", -- 0x1710
    x"60",x"C6",x"DC",x"AA",x"10",x"E0",x"85",x"D1", -- 0x1718
    x"20",x"F0",x"D0",x"A6",x"DC",x"E8",x"D0",x"02", -- 0x1720
    x"E6",x"DD",x"8A",x"48",x"46",x"DD",x"6A",x"AC", -- 0x1728
    x"61",x"03",x"C0",x"03",x"F0",x"05",x"90",x"06", -- 0x1730
    x"46",x"DD",x"6A",x"46",x"DD",x"4A",x"AC",x"1A", -- 0x1738
    x"03",x"AA",x"F0",x"0F",x"98",x"38",x"E9",x"08", -- 0x1740
    x"A8",x"B0",x"02",x"C6",x"D7",x"20",x"04",x"D1", -- 0x1748
    x"CA",x"D0",x"F1",x"68",x"2D",x"61",x"03",x"F0", -- 0x1750
    x"B5",x"AA",x"A9",x"00",x"0A",x"0D",x"63",x"03", -- 0x1758
    x"CA",x"D0",x"F9",x"85",x"D1",x"98",x"38",x"E9", -- 0x1760
    x"08",x"A8",x"B0",x"02",x"C6",x"D7",x"20",x"F3", -- 0x1768
    x"D0",x"4C",x"0E",x"D7",x"FE",x"08",x"03",x"D0", -- 0x1770
    x"03",x"FE",x"09",x"03",x"38",x"BD",x"00",x"03", -- 0x1778
    x"FD",x"02",x"03",x"9D",x"00",x"03",x"BD",x"01", -- 0x1780
    x"03",x"FD",x"03",x"03",x"9D",x"01",x"03",x"10", -- 0x1788
    x"30",x"BD",x"0A",x"03",x"30",x"0B",x"FE",x"06", -- 0x1790
    x"03",x"D0",x"11",x"FE",x"07",x"03",x"4C",x"AC", -- 0x1798
    x"D7",x"BD",x"06",x"03",x"D0",x"03",x"DE",x"07", -- 0x17A0
    x"03",x"DE",x"06",x"03",x"18",x"BD",x"00",x"03", -- 0x17A8
    x"7D",x"04",x"03",x"9D",x"00",x"03",x"BD",x"01", -- 0x17B0
    x"03",x"7D",x"05",x"03",x"9D",x"01",x"03",x"30", -- 0x17B8
    x"D0",x"60",x"AC",x"60",x"03",x"D0",x"15",x"B1", -- 0x17C0
    x"D8",x"A0",x"02",x"D9",x"B7",x"C4",x"D0",x"04", -- 0x17C8
    x"B9",x"B6",x"C4",x"88",x"88",x"10",x"F4",x"AC", -- 0x17D0
    x"55",x"03",x"AA",x"60",x"20",x"08",x"D8",x"A2", -- 0x17D8
    x"20",x"8A",x"48",x"20",x"3E",x"D0",x"68",x"AA", -- 0x17E0
    x"A0",x"07",x"B9",x"28",x"03",x"D1",x"DE",x"D0", -- 0x17E8
    x"08",x"88",x"10",x"F6",x"8A",x"E0",x"7F",x"D0", -- 0x17F0
    x"DE",x"E8",x"A5",x"DE",x"18",x"69",x"08",x"85", -- 0x17F8
    x"DE",x"D0",x"E5",x"8A",x"D0",x"DB",x"F0",x"CF", -- 0x1800
    x"A0",x"07",x"84",x"DA",x"A9",x"01",x"85",x"DB", -- 0x1808
    x"AD",x"62",x"03",x"85",x"DC",x"B1",x"D8",x"4D", -- 0x1810
    x"58",x"03",x"18",x"24",x"DC",x"F0",x"01",x"38", -- 0x1818
    x"26",x"DB",x"B0",x"0A",x"46",x"DC",x"90",x"F3", -- 0x1820
    x"98",x"69",x"07",x"A8",x"90",x"E2",x"A4",x"DA", -- 0x1828
    x"A5",x"DB",x"99",x"28",x"03",x"88",x"10",x"D2", -- 0x1830
    x"60",x"48",x"AA",x"20",x"49",x"D1",x"68",x"AA", -- 0x1838
    x"20",x"5F",x"D8",x"D0",x"15",x"B1",x"D6",x"0A", -- 0x1840
    x"26",x"DA",x"06",x"D1",x"08",x"B0",x"02",x"46", -- 0x1848
    x"DA",x"28",x"D0",x"F3",x"A5",x"DA",x"2D",x"60", -- 0x1850
    x"03",x"60",x"A9",x"FF",x"60",x"A2",x"20",x"20", -- 0x1858
    x"0F",x"D1",x"D0",x"F8",x"BD",x"02",x"03",x"49", -- 0x1860
    x"FF",x"A8",x"29",x"07",x"8D",x"1A",x"03",x"98", -- 0x1868
    x"4A",x"4A",x"4A",x"0A",x"A8",x"B1",x"E0",x"85", -- 0x1870
    x"DA",x"C8",x"B1",x"E0",x"AC",x"56",x"03",x"F0", -- 0x1878
    x"03",x"46",x"DA",x"6A",x"6D",x"50",x"03",x"85", -- 0x1880
    x"D6",x"A5",x"DA",x"6D",x"51",x"03",x"85",x"D7", -- 0x1888
    x"BD",x"01",x"03",x"85",x"DA",x"BD",x"00",x"03", -- 0x1890
    x"48",x"2D",x"61",x"03",x"6D",x"61",x"03",x"A8", -- 0x1898
    x"B9",x"06",x"C4",x"85",x"D1",x"68",x"AC",x"61", -- 0x18A0
    x"03",x"C0",x"03",x"F0",x"05",x"B0",x"06",x"0A", -- 0x18A8
    x"26",x"DA",x"0A",x"26",x"DA",x"29",x"F8",x"18", -- 0x18B0
    x"65",x"D6",x"85",x"D6",x"A5",x"DA",x"65",x"D7", -- 0x18B8
    x"10",x"04",x"38",x"ED",x"54",x"03",x"85",x"D7", -- 0x18C0
    x"AC",x"1A",x"03",x"A9",x"00",x"60",x"48",x"A9", -- 0x18C8
    x"A0",x"AE",x"6A",x"02",x"D0",x"40",x"24",x"D0", -- 0x18D0
    x"D0",x"3C",x"70",x"19",x"AD",x"5F",x"03",x"29", -- 0x18D8
    x"9F",x"09",x"40",x"20",x"54",x"C9",x"A2",x"18", -- 0x18E0
    x"A0",x"64",x"20",x"82",x"D4",x"20",x"7A",x"CD", -- 0x18E8
    x"A9",x"02",x"20",x"9D",x"C5",x"A9",x"BF",x"20", -- 0x18F0
    x"A8",x"C5",x"68",x"29",x"7F",x"20",x"C0",x"C4", -- 0x18F8
    x"A9",x"40",x"4C",x"9D",x"C5",x"A9",x"20",x"24", -- 0x1900
    x"D0",x"50",x"C0",x"D0",x"BE",x"20",x"C2",x"D7", -- 0x1908
    x"F0",x"05",x"48",x"20",x"64",x"C6",x"68",x"60", -- 0x1910
    x"A9",x"BD",x"20",x"A8",x"C5",x"20",x"51",x"C9", -- 0x1918
    x"A9",x"0D",x"60",x"AE",x"55",x"03",x"8A",x"29", -- 0x1920
    x"07",x"A8",x"BE",x"40",x"C4",x"BD",x"5E",x"C4", -- 0x1928
    x"A2",x"00",x"2C",x"8E",x"02",x"30",x"07",x"29", -- 0x1930
    x"3F",x"C0",x"04",x"B0",x"01",x"8A",x"A8",x"60", -- 0x1938
    x"10",x"E3",x"54",x"DC",x"93",x"DC",x"89",x"DE", -- 0x1940
    x"89",x"DF",x"72",x"E7",x"EB",x"E7",x"A4",x"E0", -- 0x1948
    x"C5",x"DE",x"7D",x"F2",x"8E",x"F1",x"C9",x"F4", -- 0x1950
    x"29",x"F5",x"A6",x"FF",x"CA",x"F3",x"B1",x"F1", -- 0x1958
    x"A6",x"FF",x"A6",x"FF",x"A6",x"FF",x"A6",x"FF", -- 0x1960
    x"02",x"EF",x"B3",x"E4",x"64",x"E4",x"D1",x"E1", -- 0x1968
    x"A6",x"FF",x"A6",x"FF",x"A6",x"FF",x"90",x"01", -- 0x1970
    x"9F",x"0D",x"A1",x"02",x"2B",x"F0",x"00",x"03", -- 0x1978
    x"00",x"00",x"FF",x"00",x"00",x"01",x"00",x"00", -- 0x1980
    x"00",x"00",x"00",x"FF",x"04",x"04",x"00",x"FF", -- 0x1988
    x"56",x"19",x"19",x"19",x"32",x"08",x"00",x"00", -- 0x1990
    x"00",x"00",x"20",x"09",x"00",x"00",x"00",x"00", -- 0x1998
    x"00",x"50",x"00",x"03",x"90",x"64",x"06",x"81", -- 0x19A0
    x"00",x"00",x"00",x"09",x"1B",x"01",x"D0",x"E0", -- 0x19A8
    x"F0",x"01",x"80",x"90",x"00",x"00",x"00",x"FF", -- 0x19B0
    x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x19B8
    x"00",x"00",x"64",x"05",x"FF",x"01",x"0A",x"00", -- 0x19C0
    x"00",x"00",x"00",x"00",x"FF",x"A9",x"40",x"8D", -- 0x19C8
    x"00",x"0D",x"78",x"D8",x"A2",x"FF",x"9A",x"AD", -- 0x19D0
    x"4E",x"FE",x"0A",x"48",x"F0",x"09",x"AD",x"58", -- 0x19D8
    x"02",x"4A",x"C9",x"01",x"D0",x"1D",x"4A",x"A2", -- 0x19E0
    x"04",x"86",x"01",x"85",x"00",x"A8",x"91",x"00", -- 0x19E8
    x"C5",x"01",x"F0",x"09",x"C8",x"D0",x"F7",x"C8", -- 0x19F0
    x"E8",x"E6",x"01",x"10",x"F1",x"8E",x"8E",x"02", -- 0x19F8
    x"8E",x"84",x"02",x"A2",x"0F",x"8E",x"42",x"FE", -- 0x1A00
    x"CA",x"8E",x"40",x"FE",x"E0",x"09",x"B0",x"F8", -- 0x1A08
    x"E8",x"8A",x"20",x"2A",x"F0",x"E0",x"80",x"66", -- 0x1A10
    x"FC",x"AA",x"CA",x"D0",x"F4",x"8E",x"8D",x"02", -- 0x1A18
    x"26",x"FC",x"20",x"EB",x"EE",x"6A",x"A2",x"9C", -- 0x1A20
    x"A0",x"8D",x"68",x"F0",x"09",x"A0",x"7E",x"90", -- 0x1A28
    x"11",x"A0",x"87",x"EE",x"8D",x"02",x"EE",x"8D", -- 0x1A30
    x"02",x"A5",x"FC",x"49",x"FF",x"8D",x"8F",x"02", -- 0x1A38
    x"A2",x"90",x"A9",x"00",x"E0",x"CE",x"90",x"02", -- 0x1A40
    x"A9",x"FF",x"9D",x"00",x"02",x"E8",x"D0",x"F4", -- 0x1A48
    x"8D",x"63",x"FE",x"8A",x"A2",x"E2",x"95",x"00", -- 0x1A50
    x"E8",x"D0",x"FB",x"B9",x"3F",x"D9",x"99",x"FF", -- 0x1A58
    x"01",x"88",x"D0",x"F7",x"A9",x"62",x"85",x"ED", -- 0x1A60
    x"20",x"0A",x"FB",x"A9",x"7F",x"E8",x"9D",x"4D", -- 0x1A68
    x"FE",x"9D",x"6D",x"FE",x"CA",x"10",x"F7",x"58", -- 0x1A70
    x"78",x"24",x"FC",x"50",x"03",x"20",x"55",x"F0", -- 0x1A78
    x"A2",x"F2",x"8E",x"4E",x"FE",x"A2",x"04",x"8E", -- 0x1A80
    x"4C",x"FE",x"A9",x"60",x"8D",x"4B",x"FE",x"A9", -- 0x1A88
    x"0E",x"8D",x"46",x"FE",x"8D",x"6C",x"FE",x"8D", -- 0x1A90
    x"C0",x"FE",x"CD",x"6C",x"FE",x"F0",x"03",x"EE", -- 0x1A98
    x"77",x"02",x"A9",x"27",x"8D",x"47",x"FE",x"8D", -- 0x1AA0
    x"45",x"FE",x"20",x"60",x"EC",x"AD",x"82",x"02", -- 0x1AA8
    x"29",x"7F",x"20",x"A7",x"E6",x"AE",x"84",x"02", -- 0x1AB0
    x"F0",x"03",x"20",x"C8",x"E9",x"20",x"16",x"DC", -- 0x1AB8
    x"A2",x"03",x"AC",x"07",x"80",x"B9",x"00",x"80", -- 0x1AC0
    x"DD",x"0C",x"DF",x"D0",x"2E",x"C8",x"CA",x"10", -- 0x1AC8
    x"F4",x"A6",x"F4",x"A4",x"F4",x"C8",x"C0",x"10", -- 0x1AD0
    x"B0",x"25",x"98",x"49",x"FF",x"85",x"FA",x"A9", -- 0x1AD8
    x"7F",x"85",x"FB",x"8C",x"30",x"FE",x"B1",x"FA", -- 0x1AE0
    x"8E",x"30",x"FE",x"D1",x"FA",x"D0",x"E6",x"E6", -- 0x1AE8
    x"FA",x"D0",x"F0",x"E6",x"FB",x"A5",x"FB",x"C9", -- 0x1AF0
    x"84",x"90",x"E8",x"A6",x"F4",x"10",x"0D",x"AD", -- 0x1AF8
    x"06",x"80",x"9D",x"A1",x"02",x"29",x"8F",x"D0", -- 0x1B00
    x"03",x"8E",x"4B",x"02",x"E8",x"E0",x"10",x"90", -- 0x1B08
    x"AC",x"2C",x"40",x"FE",x"30",x"11",x"CE",x"7B", -- 0x1B10
    x"02",x"A0",x"FF",x"20",x"7F",x"EE",x"CA",x"D0", -- 0x1B18
    x"F8",x"8E",x"48",x"FE",x"8E",x"49",x"FE",x"AD", -- 0x1B20
    x"8F",x"02",x"20",x"00",x"C3",x"A0",x"CA",x"20", -- 0x1B28
    x"F1",x"E4",x"20",x"D9",x"EA",x"20",x"40",x"F1", -- 0x1B30
    x"A9",x"81",x"8D",x"E0",x"FE",x"AD",x"E0",x"FE", -- 0x1B38
    x"6A",x"90",x"0A",x"A2",x"FF",x"20",x"68",x"F1", -- 0x1B40
    x"D0",x"03",x"CE",x"7A",x"02",x"A0",x"0E",x"A2", -- 0x1B48
    x"01",x"20",x"68",x"F1",x"A2",x"02",x"20",x"68", -- 0x1B50
    x"F1",x"8C",x"43",x"02",x"8C",x"44",x"02",x"A2", -- 0x1B58
    x"FE",x"AC",x"7A",x"02",x"20",x"68",x"F1",x"2D", -- 0x1B60
    x"67",x"02",x"10",x"1B",x"A0",x"02",x"20",x"A9", -- 0x1B68
    x"DE",x"AD",x"8D",x"02",x"F0",x"0C",x"A0",x"16", -- 0x1B70
    x"2C",x"8E",x"02",x"30",x"02",x"A0",x"11",x"20", -- 0x1B78
    x"A9",x"DE",x"A0",x"1B",x"20",x"A9",x"DE",x"38", -- 0x1B80
    x"20",x"D9",x"EA",x"20",x"D9",x"E9",x"08",x"68", -- 0x1B88
    x"4A",x"4A",x"4A",x"4A",x"4D",x"8F",x"02",x"29", -- 0x1B90
    x"08",x"A8",x"A2",x"03",x"20",x"68",x"F1",x"F0", -- 0x1B98
    x"1D",x"98",x"D0",x"14",x"A9",x"8D",x"20",x"35", -- 0x1BA0
    x"F1",x"A2",x"D2",x"A0",x"EA",x"CE",x"67",x"02", -- 0x1BA8
    x"20",x"F7",x"FF",x"EE",x"67",x"02",x"D0",x"06", -- 0x1BB0
    x"A9",x"00",x"AA",x"20",x"37",x"F1",x"AD",x"8D", -- 0x1BB8
    x"02",x"D0",x"05",x"AE",x"8C",x"02",x"10",x"1E", -- 0x1BC0
    x"A2",x"0F",x"BD",x"A1",x"02",x"2A",x"30",x"16", -- 0x1BC8
    x"CA",x"10",x"F7",x"A9",x"00",x"2C",x"7A",x"02", -- 0x1BD0
    x"30",x"2E",x"00",x"F9",x"4C",x"61",x"6E",x"67", -- 0x1BD8
    x"75",x"61",x"67",x"65",x"3F",x"00",x"18",x"08", -- 0x1BE0
    x"8E",x"8C",x"02",x"20",x"16",x"DC",x"A9",x"80", -- 0x1BE8
    x"A0",x"08",x"20",x"AB",x"DE",x"84",x"FD",x"20", -- 0x1BF0
    x"E7",x"FF",x"20",x"E7",x"FF",x"28",x"A9",x"01", -- 0x1BF8
    x"2C",x"7A",x"02",x"30",x"03",x"4C",x"00",x"80", -- 0x1C00
    x"4C",x"00",x"04",x"A6",x"F4",x"84",x"F4",x"8C", -- 0x1C08
    x"30",x"FE",x"A0",x"00",x"B1",x"F6",x"86",x"F4", -- 0x1C10
    x"8E",x"30",x"FE",x"60",x"85",x"FC",x"68",x"48", -- 0x1C18
    x"29",x"10",x"D0",x"03",x"6C",x"04",x"02",x"8A", -- 0x1C20
    x"48",x"BA",x"BD",x"03",x"01",x"D8",x"38",x"E9", -- 0x1C28
    x"01",x"85",x"FD",x"BD",x"04",x"01",x"E9",x"00", -- 0x1C30
    x"85",x"FE",x"A5",x"F4",x"8D",x"4A",x"02",x"86", -- 0x1C38
    x"F0",x"A2",x"06",x"20",x"68",x"F1",x"AE",x"8C", -- 0x1C40
    x"02",x"20",x"16",x"DC",x"68",x"AA",x"A5",x"FC", -- 0x1C48
    x"58",x"6C",x"02",x"02",x"A0",x"00",x"20",x"B1", -- 0x1C50
    x"DE",x"AD",x"67",x"02",x"6A",x"B0",x"FE",x"20", -- 0x1C58
    x"E7",x"FF",x"20",x"E7",x"FF",x"4C",x"B8",x"DB", -- 0x1C60
    x"38",x"6E",x"4F",x"02",x"2C",x"50",x"02",x"10", -- 0x1C68
    x"07",x"20",x"41",x"E7",x"A2",x"00",x"B0",x"02", -- 0x1C70
    x"A2",x"40",x"4C",x"7A",x"E1",x"AC",x"09",x"FE", -- 0x1C78
    x"29",x"3A",x"D0",x"34",x"AE",x"5C",x"02",x"D0", -- 0x1C80
    x"09",x"E8",x"20",x"F3",x"E4",x"20",x"41",x"E7", -- 0x1C88
    x"90",x"E6",x"60",x"D8",x"A5",x"FC",x"48",x"8A", -- 0x1C90
    x"48",x"98",x"48",x"A9",x"DE",x"48",x"A9",x"81", -- 0x1C98
    x"48",x"B8",x"AD",x"08",x"FE",x"70",x"02",x"10", -- 0x1CA0
    x"5D",x"A6",x"EA",x"CA",x"30",x"30",x"70",x"2D", -- 0x1CA8
    x"4C",x"88",x"F5",x"AC",x"09",x"FE",x"2A",x"0A", -- 0x1CB0
    x"AA",x"98",x"A0",x"07",x"4C",x"94",x"E4",x"A2", -- 0x1CB8
    x"02",x"20",x"60",x"E4",x"90",x"10",x"AD",x"85", -- 0x1CC0
    x"02",x"C9",x"02",x"D0",x"9B",x"E8",x"20",x"60", -- 0x1CC8
    x"E4",x"6E",x"D2",x"02",x"30",x"92",x"8D",x"09", -- 0x1CD0
    x"FE",x"A9",x"E7",x"85",x"EA",x"60",x"2D",x"78", -- 0x1CD8
    x"02",x"4A",x"90",x"07",x"70",x"05",x"AC",x"50", -- 0x1CE0
    x"02",x"30",x"92",x"4A",x"6A",x"B0",x"C4",x"30", -- 0x1CE8
    x"CE",x"70",x"EA",x"A2",x"05",x"20",x"68",x"F1", -- 0x1CF0
    x"F0",x"E3",x"68",x"68",x"68",x"A8",x"68",x"AA", -- 0x1CF8
    x"68",x"85",x"FC",x"6C",x"06",x"02",x"AD",x"4D", -- 0x1D00
    x"FE",x"10",x"3C",x"2D",x"79",x"02",x"2D",x"4E", -- 0x1D08
    x"FE",x"6A",x"6A",x"90",x"54",x"CE",x"40",x"02", -- 0x1D10
    x"A5",x"EA",x"10",x"02",x"E6",x"EA",x"AD",x"51", -- 0x1D18
    x"02",x"F0",x"1A",x"CE",x"51",x"02",x"D0",x"15", -- 0x1D20
    x"AE",x"52",x"02",x"AD",x"48",x"02",x"4A",x"90", -- 0x1D28
    x"03",x"AE",x"53",x"02",x"2A",x"49",x"01",x"20", -- 0x1D30
    x"00",x"EA",x"8E",x"51",x"02",x"A0",x"04",x"20", -- 0x1D38
    x"94",x"E4",x"A9",x"02",x"4C",x"6E",x"DE",x"AD", -- 0x1D40
    x"6D",x"FE",x"10",x"A7",x"2D",x"77",x"02",x"2D", -- 0x1D48
    x"6E",x"FE",x"6A",x"6A",x"90",x"9D",x"AC",x"85", -- 0x1D50
    x"02",x"88",x"D0",x"97",x"A9",x"02",x"8D",x"6D", -- 0x1D58
    x"FE",x"8D",x"6E",x"FE",x"A2",x"03",x"4C",x"3A", -- 0x1D60
    x"E1",x"2A",x"2A",x"2A",x"2A",x"10",x"5B",x"A9", -- 0x1D68
    x"20",x"A2",x"00",x"8D",x"4D",x"FE",x"8E",x"49", -- 0x1D70
    x"FE",x"A2",x"08",x"86",x"FB",x"20",x"5B",x"E4", -- 0x1D78
    x"6E",x"D7",x"02",x"30",x"44",x"A8",x"F0",x"05", -- 0x1D80
    x"20",x"6D",x"EE",x"30",x"3C",x"20",x"60",x"E4", -- 0x1D88
    x"85",x"F5",x"20",x"60",x"E4",x"85",x"F7",x"20", -- 0x1D90
    x"60",x"E4",x"85",x"F6",x"A4",x"F5",x"F0",x"1B", -- 0x1D98
    x"10",x"16",x"24",x"F5",x"70",x"05",x"20",x"BB", -- 0x1DA0
    x"EE",x"50",x"07",x"06",x"F6",x"26",x"F7",x"20", -- 0x1DA8
    x"3B",x"EE",x"AC",x"61",x"02",x"4C",x"7F",x"EE", -- 0x1DB0
    x"20",x"7F",x"EE",x"A4",x"F6",x"20",x"7F",x"EE", -- 0x1DB8
    x"A4",x"F7",x"20",x"7F",x"EE",x"46",x"FB",x"D0", -- 0x1DC0
    x"B4",x"60",x"90",x"7B",x"A9",x"40",x"8D",x"4D", -- 0x1DC8
    x"FE",x"AD",x"83",x"02",x"AA",x"49",x"0F",x"48", -- 0x1DD0
    x"A8",x"BD",x"91",x"02",x"69",x"00",x"99",x"91", -- 0x1DD8
    x"02",x"CA",x"F0",x"03",x"88",x"D0",x"F2",x"68", -- 0x1DE0
    x"8D",x"83",x"02",x"A2",x"05",x"FE",x"9B",x"02", -- 0x1DE8
    x"D0",x"08",x"CA",x"D0",x"F8",x"A0",x"05",x"20", -- 0x1DF0
    x"94",x"E4",x"AD",x"B1",x"02",x"D0",x"08",x"AD", -- 0x1DF8
    x"B2",x"02",x"F0",x"06",x"CE",x"B2",x"02",x"CE", -- 0x1E00
    x"B1",x"02",x"2C",x"CE",x"02",x"10",x"0B",x"EE", -- 0x1E08
    x"CE",x"02",x"58",x"20",x"47",x"EB",x"78",x"CE", -- 0x1E10
    x"CE",x"02",x"2C",x"D7",x"02",x"30",x"0C",x"20", -- 0x1E18
    x"6D",x"EE",x"49",x"A0",x"C9",x"60",x"90",x"03", -- 0x1E20
    x"20",x"79",x"DD",x"2C",x"B7",x"D9",x"20",x"A2", -- 0x1E28
    x"DC",x"A5",x"EC",x"05",x"ED",x"2D",x"42",x"02", -- 0x1E30
    x"F0",x"04",x"38",x"20",x"65",x"F0",x"20",x"9B", -- 0x1E38
    x"E1",x"2C",x"C0",x"FE",x"70",x"04",x"60",x"2A", -- 0x1E40
    x"10",x"28",x"AE",x"4C",x"02",x"F0",x"1D",x"AD", -- 0x1E48
    x"C2",x"FE",x"9D",x"B5",x"02",x"AD",x"C1",x"FE", -- 0x1E50
    x"9D",x"B9",x"02",x"8E",x"BE",x"02",x"A0",x"03", -- 0x1E58
    x"20",x"94",x"E4",x"CA",x"D0",x"03",x"AE",x"4D", -- 0x1E60
    x"02",x"20",x"8F",x"DE",x"A9",x"10",x"8D",x"4D", -- 0x1E68
    x"FE",x"60",x"2A",x"2A",x"2A",x"2A",x"10",x"07", -- 0x1E70
    x"20",x"65",x"F0",x"A9",x"01",x"D0",x"EF",x"4C", -- 0x1E78
    x"F3",x"DC",x"68",x"A8",x"68",x"AA",x"68",x"85", -- 0x1E80
    x"FC",x"A5",x"FC",x"40",x"8C",x"BE",x"02",x"E0", -- 0x1E88
    x"05",x"90",x"02",x"A2",x"04",x"8E",x"4C",x"02", -- 0x1E90
    x"AC",x"4E",x"02",x"88",x"98",x"29",x"08",x"18", -- 0x1E98
    x"6D",x"4C",x"02",x"E9",x"00",x"8D",x"C0",x"FE", -- 0x1EA0
    x"60",x"A9",x"C3",x"85",x"FE",x"A9",x"00",x"85", -- 0x1EA8
    x"FD",x"C8",x"B1",x"FD",x"20",x"E3",x"FF",x"AA", -- 0x1EB0
    x"D0",x"F7",x"60",x"8E",x"B1",x"02",x"8C",x"B2", -- 0x1EB8
    x"02",x"A9",x"FF",x"D0",x"02",x"A9",x"00",x"85", -- 0x1EC0
    x"E6",x"8A",x"48",x"98",x"48",x"AC",x"56",x"02", -- 0x1EC8
    x"F0",x"14",x"38",x"66",x"EB",x"20",x"D7",x"FF", -- 0x1ED0
    x"08",x"46",x"EB",x"28",x"90",x"25",x"A9",x"00", -- 0x1ED8
    x"8D",x"56",x"02",x"20",x"CE",x"FF",x"24",x"FF", -- 0x1EE0
    x"30",x"16",x"AE",x"41",x"02",x"20",x"77",x"E5", -- 0x1EE8
    x"90",x"11",x"24",x"E6",x"50",x"F0",x"AD",x"B1", -- 0x1EF0
    x"02",x"0D",x"B2",x"02",x"D0",x"E8",x"B0",x"05", -- 0x1EF8
    x"38",x"A9",x"1B",x"85",x"E6",x"68",x"A8",x"68", -- 0x1F00
    x"AA",x"A5",x"E6",x"60",x"29",x"43",x"28",x"00", -- 0x1F08
    x"2E",x"E0",x"31",x"05",x"46",x"58",x"E3",x"42", -- 0x1F10
    x"FF",x"42",x"41",x"53",x"49",x"43",x"E0",x"18", -- 0x1F18
    x"00",x"43",x"41",x"54",x"E0",x"31",x"05",x"43", -- 0x1F20
    x"4F",x"44",x"45",x"E3",x"48",x"88",x"45",x"58", -- 0x1F28
    x"45",x"43",x"F6",x"8D",x"00",x"48",x"45",x"4C", -- 0x1F30
    x"50",x"F0",x"B9",x"FF",x"4B",x"45",x"59",x"E3", -- 0x1F38
    x"27",x"FF",x"4C",x"4F",x"41",x"44",x"E2",x"3C", -- 0x1F40
    x"00",x"4C",x"49",x"4E",x"45",x"E6",x"59",x"01", -- 0x1F48
    x"4D",x"4F",x"54",x"4F",x"52",x"E3",x"48",x"89", -- 0x1F50
    x"4F",x"50",x"54",x"E3",x"48",x"8B",x"52",x"55", -- 0x1F58
    x"4E",x"E0",x"31",x"04",x"52",x"4F",x"4D",x"E3", -- 0x1F60
    x"48",x"8D",x"53",x"41",x"56",x"45",x"E2",x"3E", -- 0x1F68
    x"00",x"53",x"50",x"4F",x"4F",x"4C",x"E2",x"81", -- 0x1F70
    x"00",x"54",x"41",x"50",x"45",x"E3",x"48",x"8C", -- 0x1F78
    x"54",x"56",x"E3",x"48",x"90",x"E0",x"31",x"03", -- 0x1F80
    x"00",x"86",x"F2",x"84",x"F3",x"A9",x"08",x"20", -- 0x1F88
    x"31",x"E0",x"A0",x"00",x"B1",x"F2",x"C9",x"0D", -- 0x1F90
    x"F0",x"04",x"C8",x"D0",x"F7",x"60",x"A0",x"FF", -- 0x1F98
    x"20",x"39",x"E0",x"F0",x"72",x"C9",x"2A",x"F0", -- 0x1FA0
    x"F7",x"20",x"3A",x"E0",x"F0",x"69",x"C9",x"7C", -- 0x1FA8
    x"F0",x"65",x"C9",x"2F",x"D0",x"08",x"C8",x"20", -- 0x1FB0
    x"09",x"E0",x"A9",x"02",x"D0",x"73",x"84",x"E6", -- 0x1FB8
    x"A2",x"00",x"F0",x"13",x"5D",x"10",x"DF",x"29", -- 0x1FC0
    x"DF",x"D0",x"17",x"C8",x"18",x"B0",x"25",x"E8", -- 0x1FC8
    x"B1",x"F2",x"20",x"E3",x"E4",x"90",x"ED",x"BD", -- 0x1FD0
    x"10",x"DF",x"30",x"16",x"B1",x"F2",x"C9",x"2E", -- 0x1FD8
    x"F0",x"04",x"18",x"A4",x"E6",x"88",x"C8",x"E8", -- 0x1FE0
    x"E8",x"BD",x"0E",x"DF",x"F0",x"33",x"10",x"F8", -- 0x1FE8
    x"30",x"DB",x"E8",x"E8",x"CA",x"CA",x"48",x"BD", -- 0x1FF0
    x"11",x"DF",x"48",x"20",x"3A",x"E0",x"18",x"08", -- 0x1FF8
    x"20",x"04",x"E0",x"40",x"BD",x"12",x"DF",x"30", -- 0x2000
    x"0E",x"98",x"BC",x"12",x"DF",x"18",x"65",x"F2", -- 0x2008
    x"AA",x"98",x"A4",x"F3",x"90",x"01",x"C8",x"60", -- 0x2010
    x"AE",x"4B",x"02",x"30",x"04",x"38",x"4C",x"E7", -- 0x2018
    x"DB",x"A4",x"E6",x"A2",x"04",x"20",x"68",x"F1", -- 0x2020
    x"F0",x"ED",x"A5",x"E6",x"20",x"0D",x"E0",x"A9", -- 0x2028
    x"03",x"6C",x"1E",x"02",x"0A",x"29",x"01",x"10", -- 0x2030
    x"F8",x"C8",x"B1",x"F2",x"C9",x"20",x"F0",x"F9", -- 0x2038
    x"C9",x"0D",x"60",x"90",x"F5",x"20",x"3A",x"E0", -- 0x2040
    x"C9",x"2C",x"D0",x"F4",x"C8",x"60",x"20",x"3A", -- 0x2048
    x"E0",x"20",x"7D",x"E0",x"90",x"37",x"85",x"E6", -- 0x2050
    x"20",x"7C",x"E0",x"90",x"19",x"AA",x"A5",x"E6", -- 0x2058
    x"0A",x"B0",x"2A",x"0A",x"B0",x"27",x"65",x"E6", -- 0x2060
    x"B0",x"23",x"0A",x"B0",x"20",x"85",x"E6",x"8A", -- 0x2068
    x"65",x"E6",x"B0",x"19",x"90",x"E0",x"A6",x"E6", -- 0x2070
    x"C9",x"0D",x"38",x"60",x"C8",x"B1",x"F2",x"C9", -- 0x2078
    x"3A",x"B0",x"0A",x"C9",x"30",x"90",x"06",x"29", -- 0x2080
    x"0F",x"60",x"20",x"45",x"E0",x"18",x"60",x"20", -- 0x2088
    x"7D",x"E0",x"B0",x"0E",x"29",x"DF",x"C9",x"47", -- 0x2090
    x"B0",x"F0",x"C9",x"41",x"90",x"EC",x"08",x"E9", -- 0x2098
    x"37",x"28",x"C8",x"60",x"48",x"8A",x"48",x"98", -- 0x20A0
    x"48",x"BA",x"BD",x"03",x"01",x"48",x"2C",x"60", -- 0x20A8
    x"02",x"10",x"08",x"A8",x"A9",x"04",x"20",x"7E", -- 0x20B0
    x"E5",x"B0",x"52",x"18",x"A9",x"02",x"2C",x"7C", -- 0x20B8
    x"02",x"D0",x"05",x"68",x"48",x"20",x"C0",x"C4", -- 0x20C0
    x"A9",x"08",x"2C",x"7C",x"02",x"D0",x"02",x"90", -- 0x20C8
    x"05",x"68",x"48",x"20",x"14",x"E1",x"AD",x"7C", -- 0x20D0
    x"02",x"6A",x"90",x"1B",x"A4",x"EA",x"88",x"10", -- 0x20D8
    x"16",x"68",x"48",x"08",x"78",x"A2",x"02",x"48", -- 0x20E0
    x"20",x"5B",x"E4",x"90",x"03",x"20",x"70",x"E1", -- 0x20E8
    x"68",x"A2",x"02",x"20",x"F8",x"E1",x"28",x"A9", -- 0x20F0
    x"10",x"2C",x"7C",x"02",x"D0",x"0F",x"AC",x"57", -- 0x20F8
    x"02",x"F0",x"0A",x"68",x"48",x"38",x"66",x"EB", -- 0x2100
    x"20",x"D4",x"FF",x"46",x"EB",x"68",x"68",x"A8", -- 0x2108
    x"68",x"AA",x"68",x"60",x"2C",x"7C",x"02",x"70", -- 0x2110
    x"20",x"CD",x"86",x"02",x"F0",x"1B",x"08",x"78", -- 0x2118
    x"AA",x"A9",x"04",x"2C",x"7C",x"02",x"D0",x"10", -- 0x2120
    x"8A",x"A2",x"03",x"20",x"F8",x"E1",x"B0",x"08", -- 0x2128
    x"2C",x"D2",x"02",x"10",x"03",x"20",x"3A",x"E1", -- 0x2130
    x"28",x"60",x"AD",x"85",x"02",x"F0",x"6E",x"C9", -- 0x2138
    x"01",x"D0",x"21",x"20",x"60",x"E4",x"6E",x"D2", -- 0x2140
    x"02",x"30",x"45",x"A0",x"82",x"8C",x"6E",x"FE", -- 0x2148
    x"8D",x"61",x"FE",x"AD",x"6C",x"FE",x"29",x"F1", -- 0x2150
    x"09",x"0C",x"8D",x"6C",x"FE",x"09",x"0E",x"8D", -- 0x2158
    x"6C",x"FE",x"D0",x"2C",x"C9",x"02",x"D0",x"29", -- 0x2160
    x"A4",x"EA",x"88",x"10",x"40",x"4E",x"D2",x"02", -- 0x2168
    x"4E",x"4F",x"02",x"20",x"41",x"E7",x"90",x"18", -- 0x2170
    x"A2",x"20",x"A0",x"9F",x"08",x"78",x"98",x"86", -- 0x2178
    x"FA",x"2D",x"50",x"02",x"45",x"FA",x"AE",x"50", -- 0x2180
    x"02",x"8D",x"50",x"02",x"8D",x"08",x"FE",x"28", -- 0x2188
    x"60",x"18",x"A9",x"01",x"20",x"A2",x"E1",x"6E", -- 0x2190
    x"D2",x"02",x"60",x"2C",x"D2",x"02",x"30",x"FA", -- 0x2198
    x"A9",x"00",x"A2",x"03",x"AC",x"85",x"02",x"20", -- 0x21A0
    x"7E",x"E5",x"6C",x"22",x"02",x"18",x"48",x"08", -- 0x21A8
    x"78",x"B0",x"08",x"BD",x"AD",x"E9",x"10",x"03", -- 0x21B0
    x"20",x"A2",x"EC",x"38",x"7E",x"CF",x"02",x"E0", -- 0x21B8
    x"02",x"B0",x"08",x"A9",x"00",x"8D",x"68",x"02", -- 0x21C0
    x"8D",x"6A",x"02",x"20",x"3B",x"E7",x"28",x"68", -- 0x21C8
    x"60",x"50",x"07",x"BD",x"D8",x"02",x"9D",x"E1", -- 0x21D0
    x"02",x"60",x"08",x"78",x"08",x"38",x"BD",x"E1", -- 0x21D8
    x"02",x"FD",x"D8",x"02",x"B0",x"04",x"38",x"FD", -- 0x21E0
    x"47",x"E4",x"28",x"90",x"06",x"18",x"7D",x"47", -- 0x21E8
    x"E4",x"49",x"FF",x"A0",x"00",x"AA",x"28",x"60", -- 0x21F0
    x"78",x"20",x"B0",x"E4",x"90",x"0F",x"20",x"EA", -- 0x21F8
    x"E9",x"08",x"48",x"20",x"EB",x"EE",x"68",x"28", -- 0x2200
    x"30",x"03",x"58",x"B0",x"EB",x"60",x"48",x"A9", -- 0x2208
    x"00",x"9D",x"EE",x"02",x"9D",x"EF",x"02",x"9D", -- 0x2210
    x"F0",x"02",x"9D",x"F1",x"02",x"68",x"60",x"84", -- 0x2218
    x"E6",x"2A",x"2A",x"2A",x"2A",x"A0",x"04",x"2A", -- 0x2220
    x"3E",x"EE",x"02",x"3E",x"EF",x"02",x"3E",x"F0", -- 0x2228
    x"02",x"3E",x"F1",x"02",x"B0",x"31",x"88",x"D0", -- 0x2230
    x"EE",x"A4",x"E6",x"60",x"A9",x"FF",x"86",x"F2", -- 0x2238
    x"84",x"F3",x"8E",x"EE",x"02",x"8C",x"EF",x"02", -- 0x2240
    x"48",x"A2",x"02",x"20",x"0E",x"E2",x"A0",x"FF", -- 0x2248
    x"8C",x"F4",x"02",x"C8",x"20",x"1D",x"EA",x"20", -- 0x2250
    x"2F",x"EA",x"90",x"FB",x"68",x"48",x"F0",x"62", -- 0x2258
    x"20",x"AD",x"E2",x"B0",x"3B",x"F0",x"3E",x"00", -- 0x2260
    x"FC",x"42",x"61",x"64",x"20",x"61",x"64",x"64", -- 0x2268
    x"72",x"65",x"73",x"73",x"00",x"A2",x"10",x"20", -- 0x2270
    x"68",x"F1",x"F0",x"23",x"20",x"8B",x"F6",x"A9", -- 0x2278
    x"00",x"08",x"84",x"E6",x"AC",x"57",x"02",x"8D", -- 0x2280
    x"57",x"02",x"F0",x"03",x"20",x"CE",x"FF",x"A4", -- 0x2288
    x"E6",x"28",x"F0",x"0B",x"A9",x"80",x"20",x"CE", -- 0x2290
    x"FF",x"A8",x"F0",x"74",x"8D",x"57",x"02",x"60", -- 0x2298
    x"D0",x"6E",x"EE",x"F4",x"02",x"A2",x"EE",x"A0", -- 0x22A0
    x"02",x"68",x"4C",x"DD",x"FF",x"20",x"3A",x"E0", -- 0x22A8
    x"20",x"8F",x"E0",x"90",x"0C",x"20",x"0E",x"E2", -- 0x22B0
    x"20",x"1F",x"E2",x"20",x"8F",x"E0",x"B0",x"F8", -- 0x22B8
    x"38",x"60",x"A2",x"0A",x"20",x"AD",x"E2",x"90", -- 0x22C0
    x"47",x"B8",x"B1",x"F2",x"C9",x"2B",x"D0",x"04", -- 0x22C8
    x"2C",x"B7",x"D9",x"C8",x"A2",x"0E",x"20",x"AD", -- 0x22D0
    x"E2",x"90",x"35",x"08",x"50",x"0F",x"A2",x"FC", -- 0x22D8
    x"18",x"BD",x"FC",x"01",x"7D",x"00",x"02",x"9D", -- 0x22E0
    x"00",x"02",x"E8",x"D0",x"F4",x"A2",x"03",x"BD", -- 0x22E8
    x"F8",x"02",x"9D",x"F4",x"02",x"9D",x"F0",x"02", -- 0x22F0
    x"CA",x"10",x"F4",x"28",x"F0",x"A7",x"A2",x"06", -- 0x22F8
    x"20",x"AD",x"E2",x"90",x"0B",x"F0",x"9E",x"A2", -- 0x2300
    x"02",x"20",x"AD",x"E2",x"90",x"02",x"F0",x"95", -- 0x2308
    x"00",x"FE",x"42",x"61",x"64",x"20",x"63",x"6F", -- 0x2310
    x"6D",x"6D",x"61",x"6E",x"64",x"00",x"FB",x"42", -- 0x2318
    x"61",x"64",x"20",x"6B",x"65",x"79",x"00",x"20", -- 0x2320
    x"4E",x"E0",x"90",x"F1",x"E0",x"10",x"B0",x"ED", -- 0x2328
    x"20",x"45",x"E0",x"08",x"AE",x"10",x"0B",x"98", -- 0x2330
    x"48",x"20",x"D1",x"E3",x"68",x"A8",x"28",x"D0", -- 0x2338
    x"36",x"60",x"20",x"4E",x"E0",x"90",x"C9",x"8A", -- 0x2340
    x"48",x"A9",x"00",x"85",x"E5",x"85",x"E4",x"20", -- 0x2348
    x"43",x"E0",x"F0",x"18",x"20",x"4E",x"E0",x"90", -- 0x2350
    x"B7",x"86",x"E5",x"20",x"45",x"E0",x"F0",x"0C", -- 0x2358
    x"20",x"4E",x"E0",x"90",x"AB",x"86",x"E4",x"20", -- 0x2360
    x"3A",x"E0",x"D0",x"A4",x"A4",x"E4",x"A6",x"E5", -- 0x2368
    x"68",x"20",x"F4",x"FF",x"70",x"9A",x"60",x"38", -- 0x2370
    x"20",x"1E",x"EA",x"20",x"2F",x"EA",x"B0",x"08", -- 0x2378
    x"E8",x"F0",x"9A",x"9D",x"00",x"0B",x"90",x"F3", -- 0x2380
    x"D0",x"93",x"08",x"78",x"20",x"D1",x"E3",x"A2", -- 0x2388
    x"10",x"E4",x"E6",x"F0",x"0E",x"BD",x"00",x"0B", -- 0x2390
    x"D9",x"00",x"0B",x"D0",x"06",x"AD",x"10",x"0B", -- 0x2398
    x"9D",x"00",x"0B",x"CA",x"10",x"EB",x"28",x"60", -- 0x23A0
    x"08",x"78",x"AD",x"10",x"0B",x"38",x"F9",x"00", -- 0x23A8
    x"0B",x"85",x"FB",x"8A",x"48",x"A2",x"10",x"BD", -- 0x23B0
    x"00",x"0B",x"38",x"F9",x"00",x"0B",x"90",x"08", -- 0x23B8
    x"F0",x"06",x"C5",x"FB",x"B0",x"02",x"85",x"FB", -- 0x23C0
    x"CA",x"10",x"EC",x"68",x"AA",x"A5",x"FB",x"28", -- 0x23C8
    x"60",x"08",x"78",x"8A",x"48",x"A4",x"E6",x"20", -- 0x23D0
    x"A8",x"E3",x"B9",x"00",x"0B",x"A8",x"18",x"65", -- 0x23D8
    x"FB",x"AA",x"85",x"FA",x"AD",x"68",x"02",x"F0", -- 0x23E0
    x"0D",x"00",x"FA",x"4B",x"65",x"79",x"20",x"69", -- 0x23E8
    x"6E",x"20",x"75",x"73",x"65",x"00",x"CE",x"84", -- 0x23F0
    x"02",x"68",x"38",x"E5",x"FA",x"85",x"FA",x"F0", -- 0x23F8
    x"0C",x"BD",x"01",x"0B",x"99",x"01",x"0B",x"C8", -- 0x2400
    x"E8",x"C6",x"FA",x"D0",x"F4",x"98",x"48",x"A4", -- 0x2408
    x"E6",x"A2",x"10",x"BD",x"00",x"0B",x"D9",x"00", -- 0x2410
    x"0B",x"90",x"07",x"F0",x"05",x"E5",x"FB",x"9D", -- 0x2418
    x"00",x"0B",x"CA",x"10",x"EE",x"AD",x"10",x"0B", -- 0x2420
    x"99",x"00",x"0B",x"68",x"8D",x"10",x"0B",x"AA", -- 0x2428
    x"EE",x"84",x"02",x"28",x"60",x"03",x"0A",x"08", -- 0x2430
    x"07",x"07",x"07",x"07",x"07",x"09",x"00",x"00", -- 0x2438
    x"C0",x"C0",x"50",x"60",x"70",x"80",x"00",x"E0", -- 0x2440
    x"00",x"40",x"C0",x"F0",x"F0",x"F0",x"F0",x"C0", -- 0x2448
    x"BD",x"3E",x"E4",x"85",x"FA",x"BD",x"35",x"E4", -- 0x2450
    x"85",x"FB",x"60",x"2C",x"B7",x"D9",x"70",x"01", -- 0x2458
    x"B8",x"6C",x"2C",x"02",x"08",x"78",x"BD",x"D8", -- 0x2460
    x"02",x"DD",x"E1",x"02",x"F0",x"72",x"A8",x"20", -- 0x2468
    x"50",x"E4",x"B1",x"FA",x"70",x"1B",x"48",x"C8", -- 0x2470
    x"98",x"D0",x"03",x"BD",x"47",x"E4",x"9D",x"D8", -- 0x2478
    x"02",x"E0",x"02",x"90",x"0A",x"DD",x"E1",x"02", -- 0x2480
    x"D0",x"05",x"A0",x"00",x"20",x"94",x"E4",x"68", -- 0x2488
    x"A8",x"28",x"18",x"60",x"08",x"78",x"48",x"85", -- 0x2490
    x"FA",x"B9",x"BF",x"02",x"F0",x"41",x"98",x"A4", -- 0x2498
    x"FA",x"20",x"A5",x"F0",x"68",x"28",x"18",x"60", -- 0x24A0
    x"98",x"A0",x"02",x"20",x"94",x"E4",x"A8",x"98", -- 0x24A8
    x"6C",x"2A",x"02",x"08",x"78",x"48",x"BC",x"E1", -- 0x24B0
    x"02",x"C8",x"D0",x"03",x"BC",x"47",x"E4",x"98", -- 0x24B8
    x"DD",x"D8",x"02",x"F0",x"0F",x"BC",x"E1",x"02", -- 0x24C0
    x"9D",x"E1",x"02",x"20",x"50",x"E4",x"68",x"91", -- 0x24C8
    x"FA",x"28",x"18",x"60",x"68",x"E0",x"02",x"B0", -- 0x24D0
    x"07",x"A0",x"01",x"20",x"94",x"E4",x"48",x"68", -- 0x24D8
    x"28",x"38",x"60",x"48",x"29",x"DF",x"C9",x"41", -- 0x24E0
    x"90",x"04",x"C9",x"5B",x"90",x"01",x"38",x"68", -- 0x24E8
    x"60",x"A2",x"00",x"8A",x"2D",x"45",x"02",x"D0", -- 0x24F0
    x"B6",x"98",x"4D",x"6C",x"02",x"0D",x"75",x"02", -- 0x24F8
    x"D0",x"A6",x"AD",x"58",x"02",x"6A",x"98",x"B0", -- 0x2500
    x"0A",x"A0",x"06",x"20",x"94",x"E4",x"90",x"03", -- 0x2508
    x"20",x"74",x"E6",x"18",x"60",x"6A",x"68",x"B0", -- 0x2510
    x"79",x"98",x"48",x"4A",x"4A",x"4A",x"4A",x"49", -- 0x2518
    x"04",x"A8",x"B9",x"65",x"02",x"C9",x"01",x"F0", -- 0x2520
    x"6B",x"68",x"90",x"0D",x"29",x"0F",x"18",x"79", -- 0x2528
    x"65",x"02",x"18",x"60",x"20",x"6F",x"E8",x"68", -- 0x2530
    x"AA",x"20",x"60",x"E4",x"B0",x"55",x"48",x"E0", -- 0x2538
    x"01",x"D0",x"06",x"20",x"73",x"E1",x"A2",x"01", -- 0x2540
    x"38",x"68",x"90",x"05",x"AC",x"45",x"02",x"D0", -- 0x2548
    x"41",x"A8",x"10",x"3E",x"29",x"0F",x"C9",x"0B", -- 0x2550
    x"90",x"BF",x"69",x"7B",x"48",x"AD",x"7D",x"02", -- 0x2558
    x"D0",x"B3",x"AD",x"7C",x"02",x"6A",x"6A",x"68", -- 0x2560
    x"B0",x"CF",x"C9",x"87",x"F0",x"38",x"A8",x"8A", -- 0x2568
    x"48",x"98",x"20",x"CE",x"D8",x"68",x"AA",x"2C", -- 0x2570
    x"5F",x"02",x"10",x"05",x"A9",x"06",x"6C",x"24", -- 0x2578
    x"02",x"AD",x"68",x"02",x"F0",x"B3",x"AC",x"C9", -- 0x2580
    x"02",x"B9",x"01",x"0B",x"EE",x"C9",x"02",x"CE", -- 0x2588
    x"68",x"02",x"18",x"60",x"68",x"29",x"0F",x"A8", -- 0x2590
    x"20",x"A8",x"E3",x"8D",x"68",x"02",x"B9",x"00", -- 0x2598
    x"0B",x"8D",x"C9",x"02",x"D0",x"D1",x"8A",x"48", -- 0x25A0
    x"20",x"05",x"D9",x"A8",x"F0",x"86",x"68",x"AA", -- 0x25A8
    x"98",x"18",x"60",x"21",x"E8",x"88",x"E9",x"D3", -- 0x25B0
    x"E6",x"97",x"E9",x"97",x"E9",x"76",x"E9",x"88", -- 0x25B8
    x"E9",x"8B",x"E6",x"89",x"E6",x"B0",x"E6",x"B2", -- 0x25C0
    x"E6",x"95",x"E9",x"8C",x"E9",x"F9",x"E6",x"FA", -- 0x25C8
    x"E6",x"A8",x"F0",x"06",x"E7",x"8C",x"DE",x"C8", -- 0x25D0
    x"E9",x"B6",x"E9",x"07",x"CD",x"B4",x"F0",x"6C", -- 0x25D8
    x"E8",x"D9",x"E9",x"75",x"E2",x"45",x"F0",x"CF", -- 0x25E0
    x"F0",x"CD",x"F0",x"97",x"E1",x"73",x"E6",x"74", -- 0x25E8
    x"E6",x"5C",x"E6",x"35",x"E0",x"4F",x"E7",x"13", -- 0x25F0
    x"E7",x"29",x"E7",x"85",x"F0",x"23",x"D9",x"26", -- 0x25F8
    x"D9",x"47",x"D6",x"C2",x"D7",x"57",x"E6",x"7F", -- 0x2600
    x"E6",x"AF",x"E4",x"34",x"E0",x"35",x"F1",x"35", -- 0x2608
    x"F1",x"E7",x"DB",x"68",x"F1",x"E3",x"EA",x"60", -- 0x2610
    x"E4",x"AA",x"FF",x"F4",x"EA",x"AE",x"FF",x"F9", -- 0x2618
    x"EA",x"B2",x"FF",x"FE",x"EA",x"5B",x"E4",x"F3", -- 0x2620
    x"E4",x"FF",x"E9",x"10",x"EA",x"7C",x"E1",x"A7", -- 0x2628
    x"FF",x"6D",x"EE",x"7F",x"EE",x"C0",x"E9",x"9C", -- 0x2630
    x"E9",x"59",x"E6",x"02",x"E9",x"D5",x"E8",x"E8", -- 0x2638
    x"E8",x"D1",x"E8",x"E4",x"E8",x"03",x"E8",x"0B", -- 0x2640
    x"E8",x"2D",x"E8",x"AE",x"E8",x"35",x"C7",x"F3", -- 0x2648
    x"CB",x"48",x"C7",x"E0",x"C8",x"CE",x"D5",x"A9", -- 0x2650
    x"00",x"6C",x"00",x"02",x"A2",x"00",x"24",x"FF", -- 0x2658
    x"10",x"11",x"AD",x"76",x"02",x"D0",x"0A",x"58", -- 0x2660
    x"8D",x"69",x"02",x"20",x"8D",x"F6",x"20",x"AA", -- 0x2668
    x"F0",x"A2",x"FF",x"18",x"66",x"FF",x"2C",x"7A", -- 0x2670
    x"02",x"30",x"01",x"60",x"4C",x"03",x"04",x"AD", -- 0x2678
    x"82",x"02",x"A8",x"2A",x"E0",x"01",x"6A",x"50", -- 0x2680
    x"1E",x"A9",x"38",x"49",x"3F",x"85",x"FA",x"AC", -- 0x2688
    x"82",x"02",x"E0",x"09",x"B0",x"17",x"3D",x"AD", -- 0x2690
    x"E9",x"85",x"FB",x"98",x"05",x"FA",x"45",x"FA", -- 0x2698
    x"05",x"FB",x"09",x"40",x"4D",x"5D",x"02",x"8D", -- 0x26A0
    x"82",x"02",x"8D",x"10",x"FE",x"98",x"AA",x"60", -- 0x26A8
    x"C8",x"18",x"B9",x"52",x"02",x"48",x"8A",x"99", -- 0x26B0
    x"52",x"02",x"68",x"A8",x"AD",x"51",x"02",x"D0", -- 0x26B8
    x"10",x"8E",x"51",x"02",x"AD",x"48",x"02",x"08", -- 0x26C0
    x"6A",x"28",x"2A",x"8D",x"48",x"02",x"8D",x"20", -- 0x26C8
    x"FE",x"50",x"DA",x"8A",x"29",x"01",x"48",x"AD", -- 0x26D0
    x"50",x"02",x"2A",x"E0",x"01",x"6A",x"CD",x"50", -- 0x26D8
    x"02",x"08",x"8D",x"50",x"02",x"8D",x"08",x"FE", -- 0x26E0
    x"20",x"73",x"E1",x"28",x"F0",x"03",x"2C",x"09", -- 0x26E8
    x"FE",x"AE",x"41",x"02",x"68",x"8D",x"41",x"02", -- 0x26F0
    x"60",x"98",x"E0",x"0A",x"B0",x"B0",x"BC",x"BF", -- 0x26F8
    x"02",x"9D",x"BF",x"02",x"50",x"A7",x"F0",x"03", -- 0x2700
    x"20",x"8C",x"DE",x"AD",x"4D",x"02",x"8E",x"4D", -- 0x2708
    x"02",x"AA",x"60",x"98",x"30",x"0B",x"58",x"20", -- 0x2710
    x"BB",x"DE",x"B0",x"03",x"AA",x"A9",x"00",x"A8", -- 0x2718
    x"60",x"8A",x"49",x"7F",x"AA",x"20",x"68",x"F0", -- 0x2720
    x"2A",x"A2",x"FF",x"A0",x"FF",x"B0",x"02",x"E8", -- 0x2728
    x"C8",x"60",x"8A",x"49",x"FF",x"AA",x"E0",x"02", -- 0x2730
    x"B8",x"50",x"03",x"2C",x"B7",x"D9",x"6C",x"2E", -- 0x2738
    x"02",x"38",x"A2",x"01",x"20",x"38",x"E7",x"C0", -- 0x2740
    x"01",x"B0",x"03",x"EC",x"5B",x"02",x"60",x"30", -- 0x2748
    x"E1",x"F0",x"0C",x"E0",x"05",x"B0",x"D2",x"BC", -- 0x2750
    x"B9",x"02",x"BD",x"B5",x"02",x"AA",x"60",x"AD", -- 0x2758
    x"40",x"FE",x"6A",x"6A",x"6A",x"6A",x"49",x"FF", -- 0x2760
    x"29",x"03",x"AC",x"BE",x"02",x"8E",x"BE",x"02", -- 0x2768
    x"AA",x"60",x"48",x"08",x"78",x"85",x"EF",x"86", -- 0x2770
    x"F0",x"84",x"F1",x"A2",x"07",x"C9",x"75",x"90", -- 0x2778
    x"41",x"C9",x"A1",x"90",x"09",x"C9",x"A6",x"90", -- 0x2780
    x"3F",x"18",x"A9",x"A1",x"69",x"00",x"38",x"E9", -- 0x2788
    x"5F",x"0A",x"38",x"84",x"F1",x"A8",x"2C",x"5E", -- 0x2790
    x"02",x"10",x"07",x"8A",x"B8",x"20",x"7E",x"E5", -- 0x2798
    x"70",x"1A",x"B9",x"B4",x"E5",x"85",x"FB",x"B9", -- 0x27A0
    x"B3",x"E5",x"85",x"FA",x"A5",x"EF",x"A4",x"F1", -- 0x27A8
    x"B0",x"04",x"A0",x"00",x"B1",x"F0",x"38",x"A6", -- 0x27B0
    x"F0",x"20",x"58",x"F0",x"6A",x"28",x"2A",x"68", -- 0x27B8
    x"B8",x"60",x"A0",x"00",x"C9",x"16",x"90",x"C9", -- 0x27C0
    x"08",x"08",x"68",x"68",x"20",x"68",x"F1",x"D0", -- 0x27C8
    x"05",x"A6",x"F0",x"4C",x"BC",x"E7",x"28",x"68", -- 0x27D0
    x"2C",x"B7",x"D9",x"60",x"A5",x"EB",x"30",x"32", -- 0x27D8
    x"A9",x"08",x"25",x"E2",x"D0",x"04",x"A9",x"88", -- 0x27E0
    x"25",x"BB",x"60",x"48",x"08",x"78",x"85",x"EF", -- 0x27E8
    x"86",x"F0",x"84",x"F1",x"A2",x"08",x"C9",x"E0", -- 0x27F0
    x"B0",x"90",x"C9",x"0E",x"B0",x"CA",x"69",x"44", -- 0x27F8
    x"0A",x"90",x"90",x"20",x"15",x"E8",x"A1",x"F9", -- 0x2800
    x"91",x"F0",x"60",x"20",x"15",x"E8",x"B1",x"F0", -- 0x2808
    x"81",x"F9",x"A9",x"00",x"60",x"85",x"FA",x"C8", -- 0x2810
    x"B1",x"F0",x"85",x"FB",x"A0",x"04",x"A2",x"01", -- 0x2818
    x"60",x"D0",x"FB",x"00",x"F7",x"4F",x"53",x"20", -- 0x2820
    x"31",x"2E",x"32",x"30",x"00",x"C8",x"B1",x"F0", -- 0x2828
    x"C9",x"FF",x"F0",x"59",x"C9",x"20",x"A2",x"08", -- 0x2830
    x"B0",x"90",x"88",x"20",x"C9",x"E8",x"09",x"04", -- 0x2838
    x"AA",x"90",x"05",x"20",x"AE",x"E1",x"A0",x"01", -- 0x2840
    x"20",x"C9",x"E8",x"85",x"FA",x"08",x"A0",x"06", -- 0x2848
    x"B1",x"F0",x"48",x"A0",x"04",x"B1",x"F0",x"48", -- 0x2850
    x"A0",x"02",x"B1",x"F0",x"2A",x"38",x"E9",x"02", -- 0x2858
    x"0A",x"0A",x"05",x"FA",x"20",x"F8",x"E1",x"90", -- 0x2860
    x"1E",x"68",x"68",x"28",x"A6",x"D0",x"60",x"08", -- 0x2868
    x"78",x"AD",x"63",x"02",x"29",x"07",x"09",x"04", -- 0x2870
    x"AA",x"AD",x"64",x"02",x"20",x"B0",x"E4",x"AD", -- 0x2878
    x"66",x"02",x"48",x"AD",x"65",x"02",x"48",x"38", -- 0x2880
    x"7E",x"00",x"08",x"30",x"17",x"08",x"C8",x"B1", -- 0x2888
    x"F0",x"48",x"C8",x"B1",x"F0",x"48",x"A0",x"00", -- 0x2890
    x"B1",x"F0",x"A2",x"08",x"20",x"F8",x"E1",x"B0", -- 0x2898
    x"C8",x"6E",x"D7",x"02",x"68",x"20",x"B0",x"E4", -- 0x28A0
    x"68",x"20",x"B0",x"E4",x"28",x"60",x"E9",x"01", -- 0x28A8
    x"0A",x"0A",x"0A",x"0A",x"09",x"0F",x"AA",x"A9", -- 0x28B0
    x"00",x"A0",x"10",x"C0",x"0E",x"B0",x"02",x"B1", -- 0x28B8
    x"F0",x"9D",x"C0",x"08",x"CA",x"88",x"D0",x"F3", -- 0x28C0
    x"60",x"B1",x"F0",x"C9",x"10",x"29",x"03",x"C8", -- 0x28C8
    x"60",x"A2",x"0F",x"D0",x"03",x"AE",x"83",x"02", -- 0x28D0
    x"A0",x"04",x"BD",x"8D",x"02",x"91",x"F0",x"E8", -- 0x28D8
    x"88",x"10",x"F7",x"60",x"A9",x"0F",x"D0",x"06", -- 0x28E0
    x"AD",x"83",x"02",x"49",x"0F",x"18",x"48",x"AA", -- 0x28E8
    x"A0",x"04",x"B1",x"F0",x"9D",x"8D",x"02",x"E8", -- 0x28F0
    x"88",x"10",x"F7",x"68",x"B0",x"E5",x"8D",x"83", -- 0x28F8
    x"02",x"60",x"A0",x"04",x"B1",x"F0",x"99",x"B1", -- 0x2900
    x"02",x"88",x"C0",x"02",x"B0",x"F6",x"B1",x"F0", -- 0x2908
    x"85",x"E9",x"88",x"8C",x"69",x"02",x"B1",x"F0", -- 0x2910
    x"85",x"E8",x"58",x"90",x"07",x"A9",x"07",x"88", -- 0x2918
    x"C8",x"20",x"EE",x"FF",x"20",x"E0",x"FF",x"B0", -- 0x2920
    x"49",x"AA",x"AD",x"7C",x"02",x"6A",x"6A",x"8A", -- 0x2928
    x"B0",x"05",x"AE",x"6A",x"02",x"D0",x"EA",x"C9", -- 0x2930
    x"7F",x"D0",x"07",x"C0",x"00",x"F0",x"E5",x"88", -- 0x2938
    x"B0",x"DF",x"C9",x"15",x"D0",x"0D",x"98",x"F0", -- 0x2940
    x"DB",x"A9",x"7F",x"20",x"EE",x"FF",x"88",x"D0", -- 0x2948
    x"FA",x"F0",x"D1",x"91",x"E8",x"C9",x"0D",x"F0", -- 0x2950
    x"13",x"CC",x"B3",x"02",x"B0",x"BF",x"CD",x"B4", -- 0x2958
    x"02",x"90",x"BC",x"CD",x"B5",x"02",x"F0",x"B8", -- 0x2960
    x"90",x"B6",x"B0",x"B3",x"20",x"E7",x"FF",x"20", -- 0x2968
    x"7E",x"E5",x"A5",x"FF",x"2A",x"60",x"58",x"78", -- 0x2970
    x"24",x"FF",x"30",x"30",x"2C",x"D2",x"02",x"10", -- 0x2978
    x"F5",x"20",x"A4",x"E1",x"A0",x"00",x"84",x"F1", -- 0x2980
    x"09",x"F0",x"D0",x"0E",x"D0",x"07",x"A2",x"32", -- 0x2988
    x"8E",x"54",x"02",x"A2",x"08",x"69",x"CF",x"18", -- 0x2990
    x"69",x"E9",x"86",x"F0",x"A8",x"B9",x"90",x"01", -- 0x2998
    x"AA",x"25",x"F1",x"45",x"F0",x"99",x"90",x"01", -- 0x29A0
    x"B9",x"91",x"01",x"A8",x"60",x"64",x"7F",x"5B", -- 0x29A8
    x"6D",x"C9",x"F6",x"D2",x"E4",x"40",x"AD",x"40", -- 0x29B0
    x"02",x"58",x"78",x"CD",x"40",x"02",x"F0",x"F9", -- 0x29B8
    x"BC",x"01",x"03",x"BD",x"00",x"03",x"AA",x"60", -- 0x29C0
    x"A9",x"10",x"8D",x"84",x"02",x"A2",x"00",x"9D", -- 0x29C8
    x"00",x"0B",x"E8",x"D0",x"FA",x"8E",x"84",x"02", -- 0x29D0
    x"60",x"08",x"78",x"A9",x"40",x"20",x"EA",x"E9", -- 0x29D8
    x"30",x"05",x"18",x"B8",x"20",x"68",x"F0",x"28", -- 0x29E0
    x"2A",x"60",x"90",x"09",x"A0",x"07",x"8C",x"40", -- 0x29E8
    x"FE",x"88",x"8C",x"40",x"FE",x"24",x"FF",x"60", -- 0x29F0
    x"08",x"78",x"8D",x"40",x"FE",x"28",x"60",x"8A", -- 0x29F8
    x"08",x"78",x"8D",x"48",x"02",x"8D",x"20",x"FE", -- 0x2A00
    x"AD",x"53",x"02",x"8D",x"51",x"02",x"28",x"60", -- 0x2A08
    x"8A",x"49",x"07",x"08",x"78",x"8D",x"49",x"02", -- 0x2A10
    x"8D",x"21",x"FE",x"28",x"60",x"18",x"66",x"E4", -- 0x2A18
    x"20",x"3A",x"E0",x"C8",x"C9",x"22",x"F0",x"02", -- 0x2A20
    x"88",x"18",x"66",x"E4",x"C9",x"0D",x"60",x"A9", -- 0x2A28
    x"00",x"85",x"E5",x"B1",x"F2",x"C9",x"0D",x"D0", -- 0x2A30
    x"06",x"24",x"E4",x"30",x"52",x"10",x"1B",x"C9", -- 0x2A38
    x"20",x"90",x"4C",x"D0",x"06",x"24",x"E4",x"30", -- 0x2A40
    x"40",x"50",x"0F",x"C9",x"22",x"D0",x"10",x"24", -- 0x2A48
    x"E4",x"10",x"36",x"C8",x"B1",x"F2",x"C9",x"22", -- 0x2A50
    x"F0",x"2F",x"20",x"3A",x"E0",x"38",x"60",x"C9", -- 0x2A58
    x"7C",x"D0",x"26",x"C8",x"B1",x"F2",x"C9",x"7C", -- 0x2A60
    x"F0",x"1F",x"C9",x"22",x"F0",x"1B",x"C9",x"21", -- 0x2A68
    x"D0",x"05",x"C8",x"A9",x"80",x"D0",x"BA",x"C9", -- 0x2A70
    x"20",x"90",x"14",x"C9",x"3F",x"F0",x"08",x"20", -- 0x2A78
    x"BF",x"EA",x"2C",x"B7",x"D9",x"70",x"03",x"A9", -- 0x2A80
    x"7F",x"B8",x"C8",x"05",x"E5",x"18",x"60",x"00", -- 0x2A88
    x"FD",x"42",x"61",x"64",x"20",x"73",x"74",x"72", -- 0x2A90
    x"69",x"6E",x"67",x"00",x"C9",x"30",x"F0",x"1E", -- 0x2A98
    x"C9",x"40",x"F0",x"1A",x"90",x"12",x"C9",x"7F", -- 0x2AA0
    x"F0",x"14",x"B0",x"10",x"49",x"30",x"C9",x"6F", -- 0x2AA8
    x"F0",x"04",x"C9",x"50",x"D0",x"02",x"49",x"1F", -- 0x2AB0
    x"C9",x"21",x"90",x"02",x"49",x"10",x"60",x"C9", -- 0x2AB8
    x"7F",x"F0",x"0E",x"B0",x"E7",x"C9",x"60",x"D0", -- 0x2AC0
    x"02",x"A9",x"5F",x"C9",x"40",x"90",x"02",x"29", -- 0x2AC8
    x"1F",x"60",x"2F",x"21",x"42",x"4F",x"4F",x"54", -- 0x2AD0
    x"0D",x"AD",x"87",x"02",x"49",x"4C",x"D0",x"13", -- 0x2AD8
    x"4C",x"87",x"02",x"AD",x"90",x"02",x"8E",x"90", -- 0x2AE0
    x"02",x"AA",x"98",x"29",x"01",x"AC",x"91",x"02", -- 0x2AE8
    x"8D",x"91",x"02",x"60",x"98",x"9D",x"00",x"FC", -- 0x2AF0
    x"60",x"98",x"9D",x"00",x"FD",x"60",x"98",x"9D", -- 0x2AF8
    x"00",x"FE",x"60",x"A9",x"04",x"9D",x"08",x"08", -- 0x2B00
    x"A9",x"C0",x"9D",x"04",x"08",x"AC",x"62",x"02", -- 0x2B08
    x"F0",x"02",x"A9",x"C0",x"38",x"E9",x"40",x"4A", -- 0x2B10
    x"4A",x"4A",x"49",x"0F",x"1D",x"3C",x"EB",x"09", -- 0x2B18
    x"10",x"08",x"78",x"A0",x"FF",x"8C",x"43",x"FE", -- 0x2B20
    x"8D",x"4F",x"FE",x"C8",x"8C",x"40",x"FE",x"A0", -- 0x2B28
    x"02",x"88",x"D0",x"FD",x"A0",x"08",x"8C",x"40", -- 0x2B30
    x"FE",x"A0",x"04",x"88",x"D0",x"FD",x"28",x"60", -- 0x2B38
    x"E0",x"C0",x"A0",x"80",x"4C",x"59",x"EC",x"A9", -- 0x2B40
    x"00",x"8D",x"3B",x"08",x"AD",x"38",x"08",x"D0", -- 0x2B48
    x"06",x"EE",x"3B",x"08",x"CE",x"38",x"08",x"A2", -- 0x2B50
    x"08",x"CA",x"BD",x"00",x"08",x"F0",x"E5",x"BD", -- 0x2B58
    x"CF",x"02",x"30",x"05",x"BD",x"18",x"08",x"D0", -- 0x2B60
    x"03",x"20",x"6B",x"EC",x"BD",x"18",x"08",x"F0", -- 0x2B68
    x"13",x"C9",x"FF",x"F0",x"12",x"DE",x"1C",x"08", -- 0x2B70
    x"D0",x"0D",x"A9",x"05",x"9D",x"1C",x"08",x"DE", -- 0x2B78
    x"18",x"08",x"D0",x"03",x"20",x"6B",x"EC",x"BD", -- 0x2B80
    x"24",x"08",x"F0",x"05",x"DE",x"24",x"08",x"D0", -- 0x2B88
    x"B3",x"BC",x"20",x"08",x"C0",x"FF",x"F0",x"AC", -- 0x2B90
    x"B9",x"C0",x"08",x"29",x"7F",x"9D",x"24",x"08", -- 0x2B98
    x"BD",x"08",x"08",x"C9",x"04",x"F0",x"60",x"BD", -- 0x2BA0
    x"08",x"08",x"18",x"7D",x"20",x"08",x"A8",x"B9", -- 0x2BA8
    x"CB",x"08",x"38",x"E9",x"3F",x"8D",x"3A",x"08", -- 0x2BB0
    x"B9",x"C7",x"08",x"8D",x"39",x"08",x"BD",x"04", -- 0x2BB8
    x"08",x"48",x"18",x"6D",x"39",x"08",x"50",x"07", -- 0x2BC0
    x"2A",x"A9",x"3F",x"B0",x"02",x"49",x"FF",x"9D", -- 0x2BC8
    x"04",x"08",x"2A",x"5D",x"04",x"08",x"10",x"09", -- 0x2BD0
    x"A9",x"3F",x"90",x"02",x"49",x"FF",x"9D",x"04", -- 0x2BD8
    x"08",x"CE",x"39",x"08",x"BD",x"04",x"08",x"38", -- 0x2BE0
    x"ED",x"3A",x"08",x"4D",x"39",x"08",x"30",x"09", -- 0x2BE8
    x"AD",x"3A",x"08",x"9D",x"04",x"08",x"FE",x"08", -- 0x2BF0
    x"08",x"68",x"5D",x"04",x"08",x"29",x"F8",x"F0", -- 0x2BF8
    x"06",x"BD",x"04",x"08",x"20",x"0A",x"EB",x"BD", -- 0x2C00
    x"10",x"08",x"C9",x"03",x"F0",x"4B",x"BD",x"14", -- 0x2C08
    x"08",x"D0",x"2A",x"FE",x"10",x"08",x"BD",x"10", -- 0x2C10
    x"08",x"C9",x"03",x"D0",x"10",x"BC",x"20",x"08", -- 0x2C18
    x"B9",x"C0",x"08",x"30",x"34",x"A9",x"00",x"9D", -- 0x2C20
    x"30",x"08",x"9D",x"10",x"08",x"BD",x"10",x"08", -- 0x2C28
    x"18",x"7D",x"20",x"08",x"A8",x"B9",x"C4",x"08", -- 0x2C30
    x"9D",x"14",x"08",x"F0",x"1C",x"DE",x"14",x"08", -- 0x2C38
    x"BD",x"20",x"08",x"18",x"7D",x"10",x"08",x"A8", -- 0x2C40
    x"B9",x"C1",x"08",x"18",x"7D",x"30",x"08",x"9D", -- 0x2C48
    x"30",x"08",x"18",x"7D",x"0C",x"08",x"20",x"01", -- 0x2C50
    x"ED",x"E0",x"04",x"F0",x"0D",x"4C",x"59",x"EB", -- 0x2C58
    x"A2",x"08",x"CA",x"20",x"A2",x"EC",x"E0",x"04", -- 0x2C60
    x"D0",x"F8",x"60",x"BD",x"08",x"08",x"C9",x"04", -- 0x2C68
    x"F0",x"05",x"A9",x"03",x"9D",x"08",x"08",x"BD", -- 0x2C70
    x"CF",x"02",x"F0",x"14",x"A9",x"00",x"9D",x"CF", -- 0x2C78
    x"02",x"A0",x"04",x"99",x"2B",x"08",x"88",x"D0", -- 0x2C80
    x"FA",x"9D",x"18",x"08",x"88",x"8C",x"38",x"08", -- 0x2C88
    x"BD",x"28",x"08",x"F0",x"46",x"AD",x"3B",x"08", -- 0x2C90
    x"F0",x"36",x"A9",x"00",x"9D",x"28",x"08",x"4C", -- 0x2C98
    x"98",x"ED",x"20",x"03",x"EB",x"98",x"9D",x"18", -- 0x2CA0
    x"08",x"9D",x"CF",x"02",x"9D",x"00",x"08",x"A0", -- 0x2CA8
    x"03",x"99",x"2C",x"08",x"88",x"10",x"FA",x"8C", -- 0x2CB0
    x"38",x"08",x"30",x"4A",x"08",x"78",x"BD",x"08", -- 0x2CB8
    x"08",x"C9",x"04",x"D0",x"0A",x"20",x"5B",x"E4", -- 0x2CC0
    x"90",x"05",x"A9",x"00",x"9D",x"00",x"08",x"28", -- 0x2CC8
    x"BC",x"20",x"08",x"C0",x"FF",x"D0",x"03",x"20", -- 0x2CD0
    x"03",x"EB",x"60",x"20",x"5B",x"E4",x"B0",x"DC", -- 0x2CD8
    x"29",x"03",x"F0",x"BB",x"AD",x"38",x"08",x"F0", -- 0x2CE0
    x"15",x"FE",x"28",x"08",x"2C",x"38",x"08",x"10", -- 0x2CE8
    x"0A",x"20",x"5B",x"E4",x"29",x"03",x"8D",x"38", -- 0x2CF0
    x"08",x"10",x"03",x"CE",x"38",x"08",x"4C",x"D0", -- 0x2CF8
    x"EC",x"DD",x"2C",x"08",x"F0",x"D4",x"9D",x"2C", -- 0x2D00
    x"08",x"E0",x"04",x"D0",x"09",x"29",x"0F",x"1D", -- 0x2D08
    x"3C",x"EB",x"08",x"4C",x"95",x"ED",x"48",x"29", -- 0x2D10
    x"03",x"8D",x"3C",x"08",x"A9",x"00",x"8D",x"3D", -- 0x2D18
    x"08",x"68",x"4A",x"4A",x"C9",x"0C",x"90",x"07", -- 0x2D20
    x"EE",x"3D",x"08",x"E9",x"0C",x"D0",x"F5",x"A8", -- 0x2D28
    x"AD",x"3D",x"08",x"48",x"B9",x"FB",x"ED",x"8D", -- 0x2D30
    x"3D",x"08",x"B9",x"07",x"EE",x"48",x"29",x"03", -- 0x2D38
    x"8D",x"3E",x"08",x"68",x"4A",x"4A",x"4A",x"4A", -- 0x2D40
    x"8D",x"3F",x"08",x"AD",x"3D",x"08",x"AC",x"3C", -- 0x2D48
    x"08",x"F0",x"0C",x"38",x"ED",x"3F",x"08",x"B0", -- 0x2D50
    x"03",x"CE",x"3E",x"08",x"88",x"D0",x"F4",x"8D", -- 0x2D58
    x"3D",x"08",x"68",x"A8",x"F0",x"09",x"4E",x"3E", -- 0x2D60
    x"08",x"6E",x"3D",x"08",x"88",x"D0",x"F7",x"AD", -- 0x2D68
    x"3D",x"08",x"18",x"7D",x"3D",x"C4",x"8D",x"3D", -- 0x2D70
    x"08",x"90",x"03",x"EE",x"3E",x"08",x"29",x"0F", -- 0x2D78
    x"1D",x"3C",x"EB",x"08",x"78",x"20",x"21",x"EB", -- 0x2D80
    x"AD",x"3D",x"08",x"4E",x"3E",x"08",x"6A",x"4E", -- 0x2D88
    x"3E",x"08",x"6A",x"4A",x"4A",x"4C",x"22",x"EB", -- 0x2D90
    x"08",x"78",x"20",x"60",x"E4",x"48",x"29",x"04", -- 0x2D98
    x"F0",x"15",x"68",x"BC",x"20",x"08",x"C0",x"FF", -- 0x2DA0
    x"D0",x"03",x"20",x"03",x"EB",x"20",x"60",x"E4", -- 0x2DA8
    x"20",x"60",x"E4",x"28",x"4C",x"F7",x"ED",x"68", -- 0x2DB0
    x"29",x"F8",x"0A",x"90",x"0B",x"49",x"FF",x"4A", -- 0x2DB8
    x"38",x"E9",x"40",x"20",x"0A",x"EB",x"A9",x"FF", -- 0x2DC0
    x"9D",x"20",x"08",x"A9",x"05",x"9D",x"1C",x"08", -- 0x2DC8
    x"A9",x"01",x"9D",x"24",x"08",x"A9",x"00",x"9D", -- 0x2DD0
    x"14",x"08",x"9D",x"08",x"08",x"9D",x"30",x"08", -- 0x2DD8
    x"A9",x"FF",x"9D",x"10",x"08",x"20",x"60",x"E4", -- 0x2DE0
    x"9D",x"0C",x"08",x"20",x"60",x"E4",x"28",x"48", -- 0x2DE8
    x"BD",x"0C",x"08",x"20",x"01",x"ED",x"68",x"9D", -- 0x2DF0
    x"18",x"08",x"60",x"F0",x"B7",x"82",x"4F",x"20", -- 0x2DF8
    x"F3",x"C8",x"A0",x"7B",x"57",x"35",x"16",x"E7", -- 0x2E00
    x"D7",x"CB",x"C3",x"B7",x"AA",x"A2",x"9A",x"92", -- 0x2E08
    x"8A",x"82",x"7A",x"A9",x"EF",x"85",x"F5",x"60", -- 0x2E10
    x"A2",x"0D",x"E6",x"F5",x"A4",x"F5",x"10",x"39", -- 0x2E18
    x"A2",x"00",x"86",x"F7",x"E8",x"86",x"F6",x"20", -- 0x2E20
    x"BB",x"EE",x"A2",x"03",x"20",x"62",x"EE",x"DD", -- 0x2E28
    x"0C",x"DF",x"D0",x"E4",x"CA",x"10",x"F5",x"A9", -- 0x2E30
    x"3E",x"85",x"F6",x"20",x"BB",x"EE",x"A2",x"FF", -- 0x2E38
    x"20",x"62",x"EE",x"A0",x"08",x"0A",x"76",x"F7", -- 0x2E40
    x"88",x"D0",x"FA",x"E8",x"F0",x"F2",x"18",x"90", -- 0x2E48
    x"6A",x"A2",x"0E",x"A4",x"F5",x"30",x"0B",x"A0", -- 0x2E50
    x"FF",x"08",x"20",x"68",x"F1",x"28",x"C9",x"01", -- 0x2E58
    x"98",x"60",x"08",x"78",x"A0",x"10",x"20",x"7F", -- 0x2E60
    x"EE",x"A0",x"00",x"F0",x"17",x"A0",x"00",x"F0", -- 0x2E68
    x"11",x"48",x"20",x"7A",x"EE",x"68",x"6A",x"6A", -- 0x2E70
    x"6A",x"6A",x"29",x"0F",x"09",x"40",x"A8",x"98", -- 0x2E78
    x"A0",x"01",x"08",x"78",x"2C",x"7B",x"02",x"10", -- 0x2E80
    x"21",x"48",x"B9",x"75",x"F0",x"8D",x"43",x"FE", -- 0x2E88
    x"68",x"8D",x"4F",x"FE",x"B9",x"77",x"F0",x"8D", -- 0x2E90
    x"40",x"FE",x"2C",x"40",x"FE",x"30",x"FB",x"AD", -- 0x2E98
    x"4F",x"FE",x"48",x"B9",x"79",x"F0",x"8D",x"40", -- 0x2EA0
    x"FE",x"68",x"28",x"A8",x"60",x"AD",x"CB",x"03", -- 0x2EA8
    x"85",x"F6",x"AD",x"CC",x"03",x"85",x"F7",x"A5", -- 0x2EB0
    x"F5",x"10",x"1E",x"08",x"78",x"A5",x"F6",x"20", -- 0x2EB8
    x"71",x"EE",x"A5",x"F5",x"85",x"FA",x"A5",x"F7", -- 0x2EC0
    x"2A",x"2A",x"46",x"FA",x"6A",x"46",x"FA",x"6A", -- 0x2EC8
    x"20",x"71",x"EE",x"A5",x"FA",x"20",x"7A",x"EE", -- 0x2ED0
    x"28",x"60",x"A2",x"FF",x"A5",x"EC",x"05",x"ED", -- 0x2ED8
    x"D0",x"06",x"A9",x"81",x"8D",x"4E",x"FE",x"E8", -- 0x2EE0
    x"8E",x"42",x"02",x"08",x"AD",x"5A",x"02",x"4A", -- 0x2EE8
    x"29",x"18",x"09",x"06",x"8D",x"40",x"FE",x"4A", -- 0x2EF0
    x"09",x"07",x"8D",x"40",x"FE",x"20",x"2E",x"F1", -- 0x2EF8
    x"68",x"60",x"50",x"0A",x"A9",x"01",x"8D",x"4E", -- 0x2F00
    x"FE",x"B0",x"08",x"4C",x"0F",x"F0",x"90",x"06", -- 0x2F08
    x"4C",x"D1",x"F0",x"EE",x"42",x"02",x"AD",x"5A", -- 0x2F10
    x"02",x"29",x"B7",x"A2",x"00",x"20",x"2A",x"F0", -- 0x2F18
    x"86",x"FA",x"B8",x"10",x"05",x"2C",x"B7",x"D9", -- 0x2F20
    x"09",x"08",x"E8",x"20",x"2A",x"F0",x"90",x"BB", -- 0x2F28
    x"10",x"02",x"09",x"40",x"8D",x"5A",x"02",x"A6", -- 0x2F30
    x"EC",x"F0",x"12",x"20",x"2A",x"F0",x"30",x"10", -- 0x2F38
    x"E4",x"EC",x"86",x"EC",x"D0",x"07",x"A2",x"00", -- 0x2F40
    x"86",x"EC",x"20",x"1F",x"F0",x"4C",x"E9",x"EF", -- 0x2F48
    x"E4",x"EC",x"D0",x"EE",x"A5",x"E7",x"F0",x"23", -- 0x2F50
    x"C6",x"E7",x"D0",x"1F",x"AD",x"CA",x"02",x"85", -- 0x2F58
    x"E7",x"AD",x"55",x"02",x"8D",x"CA",x"02",x"AD", -- 0x2F60
    x"5A",x"02",x"A6",x"EC",x"E0",x"D0",x"D0",x"0E", -- 0x2F68
    x"09",x"90",x"49",x"A0",x"8D",x"5A",x"02",x"A9", -- 0x2F70
    x"00",x"85",x"E7",x"4C",x"E9",x"EF",x"E0",x"C0", -- 0x2F78
    x"D0",x"0F",x"09",x"A0",x"24",x"FA",x"10",x"04", -- 0x2F80
    x"09",x"10",x"49",x"80",x"49",x"90",x"4C",x"74", -- 0x2F88
    x"EF",x"BD",x"AB",x"EF",x"D0",x"03",x"AD",x"6B", -- 0x2F90
    x"02",x"AE",x"5A",x"02",x"86",x"FA",x"26",x"FA", -- 0x2F98
    x"10",x"07",x"A6",x"ED",x"D0",x"A4",x"20",x"BF", -- 0x2FA0
    x"EA",x"26",x"FA",x"30",x"08",x"20",x"9C",x"EA", -- 0x2FA8
    x"26",x"FA",x"4C",x"C1",x"EF",x"26",x"FA",x"30", -- 0x2FB0
    x"0D",x"20",x"E3",x"E4",x"B0",x"08",x"20",x"9C", -- 0x2FB8
    x"EA",x"AE",x"5A",x"02",x"10",x"0B",x"26",x"FA", -- 0x2FC0
    x"10",x"07",x"A6",x"ED",x"D0",x"D6",x"20",x"9C", -- 0x2FC8
    x"EA",x"CD",x"6C",x"02",x"D0",x"07",x"AE",x"75", -- 0x2FD0
    x"02",x"D0",x"02",x"86",x"E7",x"A8",x"20",x"29", -- 0x2FD8
    x"F1",x"AD",x"59",x"02",x"D0",x"03",x"20",x"F1", -- 0x2FE0
    x"E4",x"A6",x"ED",x"F0",x"0B",x"20",x"2A",x"F0", -- 0x2FE8
    x"86",x"ED",x"30",x"04",x"A2",x"00",x"86",x"ED", -- 0x2FF0
    x"A6",x"ED",x"D0",x"16",x"A0",x"EC",x"20",x"CC", -- 0x2FF8
    x"F0",x"30",x"09",x"A5",x"EC",x"85",x"ED",x"86", -- 0x3000
    x"EC",x"20",x"1F",x"F0",x"4C",x"DA",x"EE",x"20", -- 0x3008
    x"2A",x"F0",x"A5",x"EC",x"D0",x"F6",x"A0",x"ED", -- 0x3010
    x"20",x"CC",x"F0",x"30",x"EF",x"10",x"E8",x"A2", -- 0x3018
    x"01",x"86",x"E7",x"AE",x"54",x"02",x"8E",x"CA", -- 0x3020
    x"02",x"60",x"A0",x"03",x"8C",x"40",x"FE",x"A0", -- 0x3028
    x"7F",x"8C",x"43",x"FE",x"8E",x"4F",x"FE",x"AE", -- 0x3030
    x"4F",x"FE",x"60",x"71",x"33",x"34",x"35",x"84", -- 0x3038
    x"38",x"87",x"2D",x"5E",x"8C",x"84",x"EC",x"86", -- 0x3040
    x"ED",x"60",x"00",x"80",x"77",x"65",x"74",x"37", -- 0x3048
    x"69",x"39",x"30",x"5F",x"8E",x"6C",x"FE",x"FD", -- 0x3050
    x"6C",x"FA",x"00",x"31",x"32",x"64",x"72",x"36", -- 0x3058
    x"75",x"6F",x"70",x"5B",x"8F",x"2C",x"B7",x"D9", -- 0x3060
    x"6C",x"28",x"02",x"01",x"61",x"78",x"66",x"79", -- 0x3068
    x"6A",x"6B",x"40",x"3A",x"0D",x"00",x"FF",x"01", -- 0x3070
    x"02",x"09",x"0A",x"02",x"73",x"63",x"67",x"68", -- 0x3078
    x"6E",x"6C",x"3B",x"5D",x"7F",x"AC",x"44",x"02", -- 0x3080
    x"A2",x"00",x"60",x"00",x"7A",x"20",x"76",x"62", -- 0x3088
    x"6D",x"2C",x"2E",x"2F",x"8B",x"AE",x"41",x"02", -- 0x3090
    x"4C",x"AD",x"E1",x"1B",x"81",x"82",x"83",x"85", -- 0x3098
    x"86",x"88",x"89",x"5C",x"8D",x"6C",x"20",x"02", -- 0x30A0
    x"D0",x"EB",x"A2",x"08",x"58",x"78",x"20",x"B4", -- 0x30A8
    x"F0",x"CA",x"10",x"F8",x"E0",x"09",x"90",x"E0", -- 0x30B0
    x"60",x"A2",x"09",x"20",x"68",x"F1",x"20",x"4A", -- 0x30B8
    x"FA",x"0D",x"4F",x"53",x"20",x"31",x"2E",x"32", -- 0x30C0
    x"30",x"0D",x"00",x"60",x"18",x"A2",x"10",x"B0", -- 0x30C8
    x"97",x"8A",x"10",x"05",x"20",x"2A",x"F0",x"B0", -- 0x30D0
    x"55",x"08",x"90",x"02",x"A0",x"EE",x"99",x"DF", -- 0x30D8
    x"01",x"A2",x"09",x"20",x"29",x"F1",x"A9",x"7F", -- 0x30E0
    x"8D",x"43",x"FE",x"A9",x"03",x"8D",x"40",x"FE", -- 0x30E8
    x"A9",x"0F",x"8D",x"4F",x"FE",x"A9",x"01",x"8D", -- 0x30F0
    x"4D",x"FE",x"8E",x"4F",x"FE",x"2C",x"4D",x"FE", -- 0x30F8
    x"F0",x"21",x"8A",x"D9",x"DF",x"01",x"90",x"16", -- 0x3100
    x"8D",x"4F",x"FE",x"2C",x"4F",x"FE",x"10",x"0E", -- 0x3108
    x"28",x"08",x"B0",x"13",x"48",x"59",x"00",x"00", -- 0x3110
    x"0A",x"C9",x"01",x"68",x"B0",x"09",x"18",x"69", -- 0x3118
    x"10",x"10",x"E0",x"CA",x"10",x"BD",x"8A",x"AA", -- 0x3120
    x"28",x"20",x"2E",x"F1",x"58",x"78",x"A9",x"0B", -- 0x3128
    x"8D",x"40",x"FE",x"8A",x"60",x"49",x"8C",x"0A", -- 0x3130
    x"8D",x"47",x"02",x"E0",x"03",x"4C",x"4B",x"F1", -- 0x3138
    x"08",x"A9",x"A1",x"85",x"E3",x"A9",x"19",x"8D", -- 0x3140
    x"D1",x"03",x"28",x"08",x"A9",x"06",x"20",x"31", -- 0x3148
    x"E0",x"A2",x"06",x"28",x"F0",x"01",x"CA",x"86", -- 0x3150
    x"C6",x"A2",x"0E",x"BD",x"51",x"D9",x"9D",x"11", -- 0x3158
    x"02",x"CA",x"D0",x"F7",x"86",x"C2",x"A2",x"0F", -- 0x3160
    x"A5",x"F4",x"48",x"8A",x"A2",x"0F",x"FE",x"A1", -- 0x3168
    x"02",x"DE",x"A1",x"02",x"10",x"0D",x"86",x"F4", -- 0x3170
    x"8E",x"30",x"FE",x"20",x"03",x"80",x"AA",x"F0", -- 0x3178
    x"05",x"A6",x"F4",x"CA",x"10",x"E8",x"68",x"85", -- 0x3180
    x"F4",x"8D",x"30",x"FE",x"8A",x"60",x"09",x"00", -- 0x3188
    x"D0",x"10",x"C0",x"00",x"D0",x"0C",x"A5",x"C6", -- 0x3190
    x"29",x"FB",x"0D",x"47",x"02",x"0A",x"0D",x"47", -- 0x3198
    x"02",x"4A",x"60",x"4C",x"F5",x"1D",x"F6",x"04", -- 0x31A0
    x"F3",x"0F",x"E3",x"04",x"F3",x"2A",x"F3",x"74", -- 0x31A8
    x"E2",x"C9",x"07",x"B0",x"ED",x"86",x"BC",x"0A", -- 0x31B0
    x"AA",x"BD",x"A4",x"F1",x"48",x"BD",x"A3",x"F1", -- 0x31B8
    x"48",x"A6",x"BC",x"60",x"08",x"48",x"20",x"27", -- 0x31C0
    x"FB",x"AD",x"C2",x"03",x"48",x"20",x"31",x"F6", -- 0x31C8
    x"68",x"F0",x"1A",x"A2",x"03",x"A9",x"FF",x"48", -- 0x31D0
    x"BD",x"BE",x"03",x"95",x"B0",x"68",x"35",x"B0", -- 0x31D8
    x"CA",x"10",x"F4",x"C9",x"FF",x"D0",x"06",x"20", -- 0x31E0
    x"E8",x"FA",x"4C",x"67",x"E2",x"AD",x"CA",x"03", -- 0x31E8
    x"4A",x"68",x"F0",x"0E",x"90",x"13",x"20",x"F2", -- 0x31F0
    x"FA",x"00",x"D5",x"4C",x"6F",x"63",x"6B",x"65", -- 0x31F8
    x"64",x"00",x"90",x"05",x"A9",x"03",x"8D",x"58", -- 0x3200
    x"02",x"A9",x"30",x"25",x"BB",x"F0",x"04",x"A5", -- 0x3208
    x"C1",x"D0",x"0A",x"98",x"48",x"20",x"BB",x"FB", -- 0x3210
    x"68",x"A8",x"20",x"D5",x"F7",x"20",x"B4",x"F9", -- 0x3218
    x"D0",x"33",x"20",x"69",x"FB",x"2C",x"CA",x"03", -- 0x3220
    x"30",x"08",x"20",x"6A",x"F9",x"20",x"7B",x"F7", -- 0x3228
    x"D0",x"D7",x"A0",x"0A",x"A5",x"CC",x"91",x"C8", -- 0x3230
    x"C8",x"A5",x"CD",x"91",x"C8",x"A9",x"00",x"C8", -- 0x3238
    x"91",x"C8",x"C8",x"91",x"C8",x"28",x"20",x"E8", -- 0x3240
    x"FA",x"24",x"BA",x"30",x"07",x"08",x"20",x"46", -- 0x3248
    x"FA",x"0D",x"00",x"28",x"60",x"20",x"37",x"F6", -- 0x3250
    x"D0",x"AF",x"86",x"F2",x"84",x"F3",x"A0",x"00", -- 0x3258
    x"20",x"1D",x"EA",x"A2",x"00",x"20",x"2F",x"EA", -- 0x3260
    x"B0",x"0D",x"F0",x"08",x"9D",x"D2",x"03",x"E8", -- 0x3268
    x"E0",x"0B",x"D0",x"F1",x"4C",x"8F",x"EA",x"A9", -- 0x3270
    x"00",x"9D",x"D2",x"03",x"60",x"48",x"86",x"C8", -- 0x3278
    x"84",x"C9",x"A0",x"00",x"B1",x"C8",x"AA",x"C8", -- 0x3280
    x"B1",x"C8",x"A8",x"20",x"5A",x"F2",x"A0",x"02", -- 0x3288
    x"B1",x"C8",x"99",x"BC",x"03",x"99",x"AE",x"00", -- 0x3290
    x"C8",x"C0",x"0A",x"D0",x"F3",x"68",x"F0",x"07", -- 0x3298
    x"C9",x"FF",x"D0",x"B0",x"4C",x"C4",x"F1",x"8D", -- 0x32A0
    x"C6",x"03",x"8D",x"C7",x"03",x"B1",x"C8",x"99", -- 0x32A8
    x"A6",x"00",x"C8",x"C0",x"12",x"D0",x"F6",x"8A", -- 0x32B0
    x"F0",x"BA",x"20",x"27",x"FB",x"20",x"34",x"F9", -- 0x32B8
    x"A9",x"00",x"20",x"BD",x"FB",x"20",x"E2",x"FB", -- 0x32C0
    x"38",x"A2",x"FD",x"BD",x"B7",x"FF",x"FD",x"B3", -- 0x32C8
    x"FF",x"9D",x"CB",x"02",x"E8",x"D0",x"F4",x"A8", -- 0x32D0
    x"D0",x"0E",x"EC",x"C8",x"03",x"A9",x"01",x"ED", -- 0x32D8
    x"C9",x"03",x"90",x"04",x"A2",x"80",x"D0",x"08", -- 0x32E0
    x"A9",x"01",x"8D",x"C9",x"03",x"8E",x"C8",x"03", -- 0x32E8
    x"8E",x"CA",x"03",x"20",x"EC",x"F7",x"30",x"49", -- 0x32F0
    x"20",x"6A",x"F9",x"EE",x"C6",x"03",x"D0",x"C8", -- 0x32F8
    x"EE",x"C7",x"03",x"D0",x"C3",x"20",x"5A",x"F2", -- 0x3300
    x"A2",x"FF",x"8E",x"C2",x"03",x"20",x"C4",x"F1", -- 0x3308
    x"2C",x"7A",x"02",x"10",x"0A",x"AD",x"C4",x"03", -- 0x3310
    x"2D",x"C5",x"03",x"C9",x"FF",x"D0",x"03",x"6C", -- 0x3318
    x"C2",x"03",x"A2",x"C2",x"A0",x"03",x"A9",x"04", -- 0x3320
    x"4C",x"C7",x"FB",x"A9",x"08",x"20",x"44",x"F3", -- 0x3328
    x"20",x"27",x"FB",x"A9",x"00",x"20",x"48",x"F3", -- 0x3330
    x"20",x"FC",x"FA",x"A9",x"F7",x"25",x"E2",x"85", -- 0x3338
    x"E2",x"60",x"A9",x"40",x"05",x"E2",x"D0",x"F7", -- 0x3340
    x"48",x"AD",x"47",x"02",x"F0",x"0B",x"20",x"13", -- 0x3348
    x"EE",x"20",x"18",x"EE",x"90",x"03",x"B8",x"50", -- 0x3350
    x"41",x"20",x"7B",x"F7",x"AD",x"C6",x"03",x"85", -- 0x3358
    x"B4",x"AD",x"C7",x"03",x"85",x"B5",x"A2",x"FF", -- 0x3360
    x"8E",x"DF",x"03",x"E8",x"86",x"BA",x"F0",x"06", -- 0x3368
    x"20",x"69",x"FB",x"20",x"7B",x"F7",x"AD",x"47", -- 0x3370
    x"02",x"F0",x"02",x"50",x"1D",x"68",x"48",x"F0", -- 0x3378
    x"2D",x"20",x"72",x"FA",x"D0",x"16",x"A9",x"30", -- 0x3380
    x"25",x"BB",x"F0",x"0E",x"AD",x"C6",x"03",x"C5", -- 0x3388
    x"B6",x"D0",x"09",x"AD",x"C7",x"03",x"C5",x"B7", -- 0x3390
    x"D0",x"02",x"68",x"60",x"AD",x"47",x"02",x"F0", -- 0x3398
    x"0D",x"20",x"AD",x"EE",x"A9",x"FF",x"8D",x"C6", -- 0x33A0
    x"03",x"8D",x"C7",x"03",x"D0",x"C2",x"50",x"05", -- 0x33A8
    x"A9",x"FF",x"20",x"D7",x"F7",x"A2",x"00",x"20", -- 0x33B0
    x"D9",x"F9",x"AD",x"47",x"02",x"F0",x"04",x"24", -- 0x33B8
    x"BB",x"50",x"DE",x"2C",x"CA",x"03",x"30",x"DC", -- 0x33C0
    x"10",x"A6",x"85",x"BC",x"8A",x"48",x"98",x"48", -- 0x33C8
    x"A5",x"BC",x"D0",x"1E",x"98",x"D0",x"0C",x"20", -- 0x33D0
    x"75",x"E2",x"20",x"78",x"F4",x"46",x"E2",x"06", -- 0x33D8
    x"E2",x"90",x"0C",x"4A",x"B0",x"F7",x"4A",x"B0", -- 0x33E0
    x"03",x"4C",x"B1",x"FB",x"20",x"78",x"F4",x"4C", -- 0x33E8
    x"71",x"F4",x"20",x"5A",x"F2",x"24",x"BC",x"50", -- 0x33F0
    x"3D",x"A9",x"00",x"8D",x"9E",x"03",x"8D",x"DD", -- 0x33F8
    x"03",x"8D",x"DE",x"03",x"A9",x"3E",x"20",x"3D", -- 0x3400
    x"F3",x"20",x"1A",x"FB",x"08",x"20",x"31",x"F6", -- 0x3408
    x"20",x"B4",x"F6",x"28",x"A2",x"FF",x"E8",x"BD", -- 0x3410
    x"B2",x"03",x"9D",x"A7",x"03",x"D0",x"F7",x"A9", -- 0x3418
    x"01",x"20",x"44",x"F3",x"AD",x"EA",x"02",x"0D", -- 0x3420
    x"EB",x"02",x"D0",x"03",x"20",x"42",x"F3",x"A9", -- 0x3428
    x"01",x"0D",x"47",x"02",x"D0",x"39",x"8A",x"D0", -- 0x3430
    x"03",x"4C",x"8F",x"EA",x"A2",x"FF",x"E8",x"BD", -- 0x3438
    x"D2",x"03",x"9D",x"80",x"03",x"D0",x"F7",x"A9", -- 0x3440
    x"FF",x"A2",x"08",x"9D",x"8B",x"03",x"CA",x"D0", -- 0x3448
    x"FA",x"8A",x"A2",x"14",x"9D",x"80",x"03",x"E8", -- 0x3450
    x"E0",x"1E",x"D0",x"F8",x"2E",x"97",x"03",x"20", -- 0x3458
    x"27",x"FB",x"20",x"34",x"F9",x"20",x"F2",x"FA", -- 0x3460
    x"A9",x"02",x"20",x"44",x"F3",x"A9",x"02",x"85", -- 0x3468
    x"BC",x"68",x"A8",x"68",x"AA",x"A5",x"BC",x"60", -- 0x3470
    x"A9",x"02",x"25",x"E2",x"F0",x"F9",x"A9",x"00", -- 0x3478
    x"8D",x"97",x"03",x"A9",x"80",x"AE",x"9D",x"03", -- 0x3480
    x"8E",x"96",x"03",x"8D",x"98",x"03",x"20",x"96", -- 0x3488
    x"F4",x"A9",x"FD",x"4C",x"3D",x"F3",x"20",x"1A", -- 0x3490
    x"FB",x"A2",x"11",x"BD",x"8C",x"03",x"9D",x"BE", -- 0x3498
    x"03",x"CA",x"10",x"F7",x"86",x"B2",x"86",x"B3", -- 0x34A0
    x"E8",x"86",x"B0",x"A9",x"09",x"85",x"B1",x"A2", -- 0x34A8
    x"7F",x"20",x"81",x"FB",x"8D",x"DF",x"03",x"20", -- 0x34B0
    x"8E",x"FB",x"20",x"E2",x"FB",x"20",x"EC",x"F7", -- 0x34B8
    x"EE",x"94",x"03",x"D0",x"03",x"EE",x"95",x"03", -- 0x34C0
    x"60",x"8A",x"48",x"98",x"48",x"A9",x"01",x"20", -- 0x34C8
    x"9C",x"FB",x"A5",x"E2",x"0A",x"B0",x"4C",x"0A", -- 0x34D0
    x"90",x"09",x"A9",x"80",x"20",x"44",x"F3",x"A9", -- 0x34D8
    x"FE",x"B0",x"38",x"AE",x"9E",x"03",x"E8",x"EC", -- 0x34E0
    x"EA",x"02",x"D0",x"2A",x"2C",x"EC",x"02",x"30", -- 0x34E8
    x"22",x"AD",x"ED",x"02",x"48",x"20",x"1A",x"FB", -- 0x34F0
    x"08",x"20",x"AC",x"F6",x"28",x"68",x"85",x"BC", -- 0x34F8
    x"18",x"2C",x"EC",x"02",x"10",x"17",x"AD",x"EA", -- 0x3500
    x"02",x"0D",x"EB",x"02",x"D0",x"0F",x"20",x"42", -- 0x3508
    x"F3",x"D0",x"0A",x"20",x"42",x"F3",x"CA",x"18", -- 0x3510
    x"BD",x"00",x"0A",x"85",x"BC",x"EE",x"9E",x"03", -- 0x3518
    x"4C",x"71",x"F4",x"00",x"DF",x"45",x"4F",x"46", -- 0x3520
    x"00",x"85",x"C4",x"8A",x"48",x"98",x"48",x"A9", -- 0x3528
    x"02",x"20",x"9C",x"FB",x"AE",x"9D",x"03",x"A5", -- 0x3530
    x"C4",x"9D",x"00",x"09",x"E8",x"D0",x"06",x"20", -- 0x3538
    x"96",x"F4",x"20",x"F2",x"FA",x"EE",x"9D",x"03", -- 0x3540
    x"A5",x"C4",x"4C",x"6F",x"F4",x"8A",x"F0",x"2E", -- 0x3548
    x"E0",x"03",x"F0",x"1F",x"C0",x"03",x"B0",x"06", -- 0x3550
    x"CA",x"F0",x"06",x"CA",x"F0",x"0A",x"4C",x"10", -- 0x3558
    x"E3",x"A9",x"33",x"C8",x"C8",x"C8",x"D0",x"02", -- 0x3560
    x"A9",x"CC",x"C8",x"25",x"E3",x"19",x"81",x"F5", -- 0x3568
    x"85",x"E3",x"60",x"98",x"30",x"02",x"D0",x"02", -- 0x3570
    x"A9",x"19",x"8D",x"D1",x"03",x"60",x"A8",x"F0", -- 0x3578
    x"EC",x"A1",x"00",x"22",x"11",x"00",x"88",x"CC", -- 0x3580
    x"C6",x"C0",x"AD",x"47",x"02",x"F0",x"07",x"20", -- 0x3588
    x"51",x"EE",x"A8",x"18",x"90",x"1A",x"AD",x"08", -- 0x3590
    x"FE",x"48",x"29",x"02",x"F0",x"0B",x"A4",x"CA", -- 0x3598
    x"F0",x"07",x"68",x"A5",x"BD",x"8D",x"09",x"FE", -- 0x35A0
    x"60",x"AC",x"09",x"FE",x"68",x"4A",x"4A",x"4A", -- 0x35A8
    x"A6",x"C2",x"F0",x"69",x"CA",x"D0",x"06",x"90", -- 0x35B0
    x"64",x"A0",x"02",x"D0",x"5E",x"CA",x"D0",x"13", -- 0x35B8
    x"B0",x"5B",x"98",x"20",x"78",x"FB",x"A0",x"03", -- 0x35C0
    x"C9",x"2A",x"F0",x"4F",x"20",x"50",x"FB",x"A0", -- 0x35C8
    x"01",x"D0",x"48",x"CA",x"D0",x"0C",x"B0",x"04", -- 0x35D0
    x"84",x"BD",x"F0",x"41",x"A9",x"80",x"85",x"C0", -- 0x35D8
    x"D0",x"3B",x"CA",x"D0",x"29",x"B0",x"2F",x"98", -- 0x35E0
    x"20",x"B0",x"F7",x"A4",x"BC",x"E6",x"BC",x"24", -- 0x35E8
    x"BD",x"30",x"0D",x"20",x"D3",x"FB",x"F0",x"05", -- 0x35F0
    x"8E",x"E5",x"FE",x"D0",x"03",x"8A",x"91",x"B0", -- 0x35F8
    x"C8",x"CC",x"C8",x"03",x"D0",x"17",x"A9",x"01", -- 0x3600
    x"85",x"BC",x"A0",x"05",x"D0",x"0D",x"98",x"20", -- 0x3608
    x"B0",x"F7",x"C6",x"BC",x"10",x"07",x"20",x"46", -- 0x3610
    x"FB",x"A0",x"00",x"84",x"C2",x"60",x"48",x"98", -- 0x3618
    x"48",x"8A",x"A8",x"A9",x"03",x"20",x"9C",x"FB", -- 0x3620
    x"A5",x"E2",x"29",x"40",x"AA",x"68",x"A8",x"68", -- 0x3628
    x"60",x"A9",x"00",x"85",x"B4",x"85",x"B5",x"A5", -- 0x3630
    x"B4",x"48",x"85",x"B6",x"A5",x"B5",x"48",x"85", -- 0x3638
    x"B7",x"20",x"46",x"FA",x"53",x"65",x"61",x"72", -- 0x3640
    x"63",x"68",x"69",x"6E",x"67",x"0D",x"00",x"A9", -- 0x3648
    x"FF",x"20",x"48",x"F3",x"68",x"85",x"B5",x"68", -- 0x3650
    x"85",x"B4",x"A5",x"B6",x"05",x"B7",x"D0",x"0D", -- 0x3658
    x"85",x"B4",x"85",x"B5",x"A5",x"C1",x"D0",x"05", -- 0x3660
    x"A2",x"B1",x"20",x"81",x"FB",x"AD",x"47",x"02", -- 0x3668
    x"F0",x"13",x"70",x"11",x"00",x"D6",x"46",x"69", -- 0x3670
    x"6C",x"65",x"20",x"6E",x"6F",x"74",x"20",x"66", -- 0x3678
    x"6F",x"75",x"6E",x"64",x"00",x"A0",x"FF",x"8C", -- 0x3680
    x"DF",x"03",x"60",x"A9",x"00",x"08",x"84",x"E6", -- 0x3688
    x"AC",x"56",x"02",x"8D",x"56",x"02",x"F0",x"03", -- 0x3690
    x"20",x"CE",x"FF",x"A4",x"E6",x"28",x"F0",x"0B", -- 0x3698
    x"A9",x"40",x"20",x"CE",x"FF",x"A8",x"F0",x"CC", -- 0x36A0
    x"8D",x"56",x"02",x"60",x"A2",x"A6",x"20",x"81", -- 0x36A8
    x"FB",x"20",x"7B",x"F7",x"AD",x"CA",x"03",x"4A", -- 0x36B0
    x"90",x"03",x"4C",x"F6",x"F1",x"AD",x"DD",x"03", -- 0x36B8
    x"85",x"B4",x"AD",x"DE",x"03",x"85",x"B5",x"A9", -- 0x36C0
    x"00",x"85",x"B0",x"A9",x"0A",x"85",x"B1",x"A9", -- 0x36C8
    x"FF",x"85",x"B2",x"85",x"B3",x"20",x"D5",x"F7", -- 0x36D0
    x"20",x"B4",x"F9",x"D0",x"25",x"AD",x"FF",x"0A", -- 0x36D8
    x"8D",x"ED",x"02",x"20",x"69",x"FB",x"8E",x"DD", -- 0x36E0
    x"03",x"8C",x"DE",x"03",x"A2",x"02",x"BD",x"C8", -- 0x36E8
    x"03",x"9D",x"EA",x"02",x"CA",x"10",x"F7",x"2C", -- 0x36F0
    x"EC",x"02",x"10",x"03",x"20",x"49",x"F2",x"4C", -- 0x36F8
    x"F2",x"FA",x"20",x"37",x"F6",x"D0",x"AD",x"C9", -- 0x3700
    x"2A",x"F0",x"37",x"C9",x"23",x"D0",x"0F",x"EE", -- 0x3708
    x"C6",x"03",x"D0",x"03",x"EE",x"C7",x"03",x"A2", -- 0x3710
    x"FF",x"2C",x"B7",x"D9",x"D0",x"55",x"A9",x"F7", -- 0x3718
    x"20",x"3D",x"F3",x"00",x"D7",x"42",x"61",x"64", -- 0x3720
    x"20",x"52",x"4F",x"4D",x"00",x"A0",x"FF",x"20", -- 0x3728
    x"90",x"FB",x"A9",x"01",x"85",x"C2",x"20",x"50", -- 0x3730
    x"FB",x"20",x"95",x"F9",x"A9",x"03",x"C5",x"C2", -- 0x3738
    x"D0",x"F7",x"A0",x"00",x"20",x"7C",x"FB",x"20", -- 0x3740
    x"97",x"F7",x"50",x"1A",x"99",x"B2",x"03",x"F0", -- 0x3748
    x"06",x"C8",x"C0",x"0B",x"D0",x"F1",x"88",x"A2", -- 0x3750
    x"0C",x"20",x"97",x"F7",x"50",x"08",x"9D",x"B2", -- 0x3758
    x"03",x"E8",x"E0",x"1F",x"D0",x"F3",x"98",x"AA", -- 0x3760
    x"A9",x"00",x"99",x"B2",x"03",x"A5",x"BE",x"05", -- 0x3768
    x"BF",x"85",x"C1",x"20",x"78",x"FB",x"84",x"C2", -- 0x3770
    x"8A",x"D0",x"59",x"AD",x"47",x"02",x"F0",x"AD", -- 0x3778
    x"20",x"51",x"EE",x"C9",x"2B",x"D0",x"80",x"A9", -- 0x3780
    x"08",x"25",x"E2",x"F0",x"03",x"20",x"4D",x"F2", -- 0x3788
    x"20",x"18",x"EE",x"90",x"EB",x"B8",x"60",x"AD", -- 0x3790
    x"47",x"02",x"F0",x"11",x"8A",x"48",x"98",x"48", -- 0x3798
    x"20",x"51",x"EE",x"85",x"BD",x"A9",x"FF",x"85", -- 0x37A0
    x"C0",x"68",x"A8",x"68",x"AA",x"20",x"84",x"F8", -- 0x37A8
    x"08",x"48",x"38",x"66",x"CB",x"45",x"BF",x"85", -- 0x37B0
    x"BF",x"A5",x"BF",x"2A",x"90",x"0C",x"6A",x"49", -- 0x37B8
    x"08",x"85",x"BF",x"A5",x"BE",x"49",x"10",x"85", -- 0x37C0
    x"BE",x"38",x"26",x"BE",x"26",x"BF",x"46",x"CB", -- 0x37C8
    x"D0",x"E7",x"68",x"28",x"60",x"A9",x"00",x"85", -- 0x37D0
    x"BD",x"A2",x"00",x"86",x"BC",x"50",x"0A",x"AD", -- 0x37D8
    x"C8",x"03",x"0D",x"C9",x"03",x"F0",x"02",x"A2", -- 0x37E0
    x"04",x"86",x"C2",x"60",x"08",x"A2",x"03",x"A9", -- 0x37E8
    x"00",x"9D",x"CB",x"03",x"CA",x"10",x"FA",x"AD", -- 0x37F0
    x"C6",x"03",x"0D",x"C7",x"03",x"D0",x"05",x"20", -- 0x37F8
    x"92",x"F8",x"F0",x"03",x"20",x"96",x"F8",x"A9", -- 0x3800
    x"2A",x"85",x"BD",x"20",x"78",x"FB",x"20",x"4A", -- 0x3808
    x"FB",x"20",x"84",x"F8",x"88",x"C8",x"B9",x"D2", -- 0x3810
    x"03",x"99",x"B2",x"03",x"20",x"75",x"F8",x"D0", -- 0x3818
    x"F4",x"A2",x"0C",x"BD",x"B2",x"03",x"20",x"75", -- 0x3820
    x"F8",x"E8",x"E0",x"1D",x"D0",x"F5",x"20",x"7B", -- 0x3828
    x"F8",x"AD",x"C8",x"03",x"0D",x"C9",x"03",x"F0", -- 0x3830
    x"1C",x"A0",x"00",x"20",x"7C",x"FB",x"B1",x"B0", -- 0x3838
    x"20",x"D3",x"FB",x"F0",x"03",x"AE",x"E5",x"FE", -- 0x3840
    x"8A",x"20",x"75",x"F8",x"C8",x"CC",x"C8",x"03", -- 0x3848
    x"D0",x"EC",x"20",x"7B",x"F8",x"20",x"84",x"F8", -- 0x3850
    x"20",x"84",x"F8",x"20",x"46",x"FB",x"A9",x"01", -- 0x3858
    x"20",x"98",x"F8",x"28",x"20",x"B9",x"F8",x"2C", -- 0x3860
    x"CA",x"03",x"10",x"08",x"08",x"20",x"92",x"F8", -- 0x3868
    x"20",x"46",x"F2",x"28",x"60",x"20",x"82",x"F8", -- 0x3870
    x"4C",x"B0",x"F7",x"A5",x"BF",x"20",x"82",x"F8", -- 0x3878
    x"A5",x"BE",x"85",x"BD",x"20",x"95",x"F9",x"24", -- 0x3880
    x"C0",x"10",x"F9",x"A9",x"00",x"85",x"C0",x"A5", -- 0x3888
    x"BD",x"60",x"A9",x"32",x"D0",x"02",x"A5",x"C7", -- 0x3890
    x"A2",x"05",x"8D",x"40",x"02",x"20",x"95",x"F9", -- 0x3898
    x"2C",x"40",x"02",x"10",x"F8",x"CA",x"D0",x"F2", -- 0x38A0
    x"60",x"AD",x"C6",x"03",x"0D",x"C7",x"03",x"F0", -- 0x38A8
    x"05",x"2C",x"DF",x"03",x"10",x"03",x"20",x"49", -- 0x38B0
    x"F2",x"A0",x"00",x"84",x"BA",x"AD",x"CA",x"03", -- 0x38B8
    x"8D",x"DF",x"03",x"20",x"DC",x"E7",x"F0",x"6B", -- 0x38C0
    x"A9",x"0D",x"20",x"EE",x"FF",x"B9",x"B2",x"03", -- 0x38C8
    x"F0",x"10",x"C9",x"20",x"90",x"04",x"C9",x"7F", -- 0x38D0
    x"90",x"02",x"A9",x"3F",x"20",x"EE",x"FF",x"C8", -- 0x38D8
    x"D0",x"EB",x"AD",x"47",x"02",x"F0",x"04",x"24", -- 0x38E0
    x"BB",x"50",x"48",x"20",x"91",x"F9",x"C8",x"C0", -- 0x38E8
    x"0B",x"90",x"EF",x"AD",x"C6",x"03",x"AA",x"20", -- 0x38F0
    x"7A",x"F9",x"2C",x"CA",x"03",x"10",x"34",x"8A", -- 0x38F8
    x"18",x"6D",x"C9",x"03",x"85",x"CD",x"20",x"75", -- 0x3900
    x"F9",x"AD",x"C8",x"03",x"85",x"CC",x"20",x"7A", -- 0x3908
    x"F9",x"24",x"BB",x"50",x"1E",x"A2",x"04",x"20", -- 0x3910
    x"91",x"F9",x"CA",x"D0",x"FA",x"A2",x"0F",x"20", -- 0x3918
    x"27",x"F9",x"20",x"91",x"F9",x"A2",x"13",x"A0", -- 0x3920
    x"04",x"BD",x"B2",x"03",x"20",x"7A",x"F9",x"CA", -- 0x3928
    x"88",x"D0",x"F6",x"60",x"AD",x"47",x"02",x"F0", -- 0x3930
    x"03",x"4C",x"10",x"E3",x"20",x"8E",x"FB",x"20", -- 0x3938
    x"E2",x"FB",x"20",x"DC",x"E7",x"F0",x"EC",x"20", -- 0x3940
    x"46",x"FA",x"52",x"45",x"43",x"4F",x"52",x"44", -- 0x3948
    x"20",x"74",x"68",x"65",x"6E",x"20",x"52",x"45", -- 0x3950
    x"54",x"55",x"52",x"4E",x"00",x"20",x"95",x"F9", -- 0x3958
    x"20",x"E0",x"FF",x"C9",x"0D",x"D0",x"F6",x"4C", -- 0x3960
    x"E7",x"FF",x"E6",x"B1",x"D0",x"06",x"E6",x"B2", -- 0x3968
    x"D0",x"02",x"E6",x"B3",x"60",x"48",x"20",x"91", -- 0x3970
    x"F9",x"68",x"48",x"4A",x"4A",x"4A",x"4A",x"20", -- 0x3978
    x"83",x"F9",x"68",x"18",x"29",x"0F",x"69",x"30", -- 0x3980
    x"C9",x"3A",x"90",x"02",x"69",x"06",x"4C",x"EE", -- 0x3988
    x"FF",x"A9",x"20",x"D0",x"F9",x"08",x"24",x"EB", -- 0x3990
    x"30",x"04",x"24",x"FF",x"30",x"02",x"28",x"60", -- 0x3998
    x"20",x"3B",x"F3",x"20",x"F2",x"FA",x"A9",x"7E", -- 0x39A0
    x"20",x"F4",x"FF",x"00",x"11",x"45",x"73",x"63", -- 0x39A8
    x"61",x"70",x"65",x"00",x"98",x"F0",x"0D",x"20", -- 0x39B0
    x"46",x"FA",x"0D",x"4C",x"6F",x"61",x"64",x"69", -- 0x39B8
    x"6E",x"67",x"0D",x"00",x"85",x"BA",x"A2",x"FF", -- 0x39C0
    x"A5",x"C1",x"D0",x"0D",x"20",x"72",x"FA",x"08", -- 0x39C8
    x"A2",x"FF",x"A0",x"99",x"A9",x"FA",x"28",x"D0", -- 0x39D0
    x"1C",x"A0",x"8E",x"A5",x"C1",x"F0",x"04",x"A9", -- 0x39D8
    x"FA",x"D0",x"12",x"AD",x"C6",x"03",x"C5",x"B4", -- 0x39E0
    x"D0",x"07",x"AD",x"C7",x"03",x"C5",x"B5",x"F0", -- 0x39E8
    x"13",x"A0",x"A4",x"A9",x"FA",x"48",x"98",x"48", -- 0x39F0
    x"8A",x"48",x"20",x"B6",x"F8",x"68",x"AA",x"68", -- 0x39F8
    x"A8",x"68",x"D0",x"14",x"8A",x"48",x"20",x"A9", -- 0x3A00
    x"F8",x"20",x"D6",x"FA",x"68",x"AA",x"A5",x"BE", -- 0x3A08
    x"05",x"BF",x"F0",x"79",x"A0",x"8E",x"A9",x"FA", -- 0x3A10
    x"C6",x"BA",x"48",x"24",x"EB",x"30",x"0D",x"8A", -- 0x3A18
    x"2D",x"47",x"02",x"D0",x"07",x"8A",x"29",x"11", -- 0x3A20
    x"25",x"BB",x"F0",x"10",x"68",x"85",x"B9",x"84", -- 0x3A28
    x"B8",x"20",x"8B",x"F6",x"46",x"EB",x"20",x"E8", -- 0x3A30
    x"FA",x"6C",x"B8",x"00",x"68",x"C8",x"D0",x"03", -- 0x3A38
    x"18",x"69",x"01",x"48",x"98",x"48",x"20",x"DC", -- 0x3A40
    x"E7",x"A8",x"68",x"85",x"B8",x"68",x"85",x"B9", -- 0x3A48
    x"98",x"08",x"E6",x"B8",x"D0",x"02",x"E6",x"B9", -- 0x3A50
    x"A0",x"00",x"B1",x"B8",x"F0",x"0A",x"28",x"08", -- 0x3A58
    x"F0",x"F0",x"20",x"E3",x"FF",x"4C",x"52",x"FA", -- 0x3A60
    x"28",x"E6",x"B8",x"D0",x"02",x"E6",x"B9",x"6C", -- 0x3A68
    x"B8",x"00",x"A2",x"FF",x"E8",x"BD",x"D2",x"03", -- 0x3A70
    x"D0",x"07",x"8A",x"F0",x"03",x"BD",x"B2",x"03", -- 0x3A78
    x"60",x"20",x"E3",x"E4",x"5D",x"B2",x"03",x"B0", -- 0x3A80
    x"02",x"29",x"DF",x"F0",x"E7",x"60",x"00",x"D8", -- 0x3A88
    x"0D",x"44",x"61",x"74",x"61",x"3F",x"00",x"D0", -- 0x3A90
    x"15",x"00",x"DB",x"0D",x"46",x"69",x"6C",x"65", -- 0x3A98
    x"3F",x"00",x"D0",x"0A",x"00",x"DA",x"0D",x"42", -- 0x3AA0
    x"6C",x"6F",x"63",x"6B",x"3F",x"00",x"A5",x"BA", -- 0x3AA8
    x"F0",x"21",x"8A",x"F0",x"1E",x"A9",x"22",x"24", -- 0x3AB0
    x"BB",x"F0",x"18",x"20",x"46",x"FB",x"A8",x"20", -- 0x3AB8
    x"4A",x"FA",x"0D",x"07",x"52",x"65",x"77",x"69", -- 0x3AC0
    x"6E",x"64",x"20",x"74",x"61",x"70",x"65",x"0D", -- 0x3AC8
    x"0D",x"00",x"60",x"20",x"4D",x"F2",x"A5",x"C2", -- 0x3AD0
    x"F0",x"F8",x"20",x"95",x"F9",x"AD",x"47",x"02", -- 0x3AD8
    x"F0",x"F4",x"20",x"88",x"F5",x"4C",x"D6",x"FA", -- 0x3AE0
    x"20",x"DC",x"E7",x"F0",x"05",x"A9",x"07",x"20", -- 0x3AE8
    x"EE",x"FF",x"A9",x"80",x"20",x"BD",x"FB",x"A2", -- 0x3AF0
    x"00",x"20",x"95",x"FB",x"08",x"78",x"AD",x"82", -- 0x3AF8
    x"02",x"8D",x"10",x"FE",x"A9",x"00",x"85",x"EA", -- 0x3B00
    x"F0",x"01",x"08",x"20",x"46",x"FB",x"AD",x"50", -- 0x3B08
    x"02",x"4C",x"89",x"E1",x"28",x"24",x"FF",x"10", -- 0x3B10
    x"18",x"60",x"A5",x"E3",x"0A",x"0A",x"0A",x"0A", -- 0x3B18
    x"85",x"BB",x"AD",x"D1",x"03",x"D0",x"08",x"A5", -- 0x3B20
    x"E3",x"29",x"F0",x"85",x"BB",x"A9",x"06",x"85", -- 0x3B28
    x"C7",x"58",x"08",x"78",x"2C",x"4F",x"02",x"10", -- 0x3B30
    x"DB",x"A5",x"EA",x"30",x"D7",x"A9",x"01",x"85", -- 0x3B38
    x"EA",x"20",x"46",x"FB",x"28",x"60",x"A9",x"03", -- 0x3B40
    x"D0",x"1B",x"A9",x"30",x"85",x"CA",x"D0",x"13", -- 0x3B48
    x"A9",x"05",x"8D",x"10",x"FE",x"A2",x"FF",x"CA", -- 0x3B50
    x"D0",x"FD",x"86",x"CA",x"A9",x"85",x"8D",x"10", -- 0x3B58
    x"FE",x"A9",x"D0",x"05",x"C6",x"8D",x"08",x"FE", -- 0x3B60
    x"60",x"AE",x"C6",x"03",x"AC",x"C7",x"03",x"E8", -- 0x3B68
    x"86",x"B4",x"D0",x"01",x"C8",x"84",x"B5",x"60", -- 0x3B70
    x"A0",x"00",x"84",x"C0",x"84",x"BE",x"84",x"BF", -- 0x3B78
    x"60",x"A0",x"FF",x"C8",x"E8",x"BD",x"00",x"03", -- 0x3B80
    x"99",x"D2",x"03",x"D0",x"F6",x"60",x"A0",x"00", -- 0x3B88
    x"58",x"A2",x"01",x"84",x"C3",x"A9",x"89",x"A4", -- 0x3B90
    x"C3",x"4C",x"F4",x"FF",x"85",x"BC",x"98",x"4D", -- 0x3B98
    x"47",x"02",x"A8",x"A5",x"E2",x"25",x"BC",x"4A", -- 0x3BA0
    x"88",x"F0",x"04",x"4A",x"88",x"D0",x"02",x"B0", -- 0x3BA8
    x"4D",x"00",x"DE",x"43",x"68",x"61",x"6E",x"6E", -- 0x3BB0
    x"65",x"6C",x"00",x"A9",x"01",x"20",x"D3",x"FB", -- 0x3BB8
    x"F0",x"3C",x"8A",x"A2",x"B0",x"A0",x"00",x"48", -- 0x3BC0
    x"A9",x"C0",x"20",x"06",x"04",x"90",x"FB",x"68", -- 0x3BC8
    x"4C",x"06",x"04",x"AA",x"A5",x"B2",x"25",x"B3", -- 0x3BD0
    x"C9",x"FF",x"F0",x"05",x"AD",x"7A",x"02",x"29", -- 0x3BD8
    x"80",x"60",x"A9",x"85",x"8D",x"10",x"FE",x"20", -- 0x3BE0
    x"46",x"FB",x"A9",x"10",x"20",x"63",x"FB",x"20", -- 0x3BE8
    x"95",x"F9",x"AD",x"08",x"FE",x"29",x"02",x"F0", -- 0x3BF0
    x"F6",x"A9",x"AA",x"8D",x"09",x"FE",x"60",x"00", -- 0x3BF8
    x"28",x"43",x"29",x"20",x"31",x"39",x"38",x"31", -- 0x3C00
    x"20",x"41",x"63",x"6F",x"72",x"6E",x"20",x"43", -- 0x3C08
    x"6F",x"6D",x"70",x"75",x"74",x"65",x"72",x"73", -- 0x3C10
    x"20",x"4C",x"74",x"64",x"2E",x"54",x"68",x"61", -- 0x3C18
    x"6E",x"6B",x"73",x"20",x"61",x"72",x"65",x"20", -- 0x3C20
    x"64",x"75",x"65",x"20",x"74",x"6F",x"20",x"74", -- 0x3C28
    x"68",x"65",x"20",x"66",x"6F",x"6C",x"6C",x"6F", -- 0x3C30
    x"77",x"69",x"6E",x"67",x"20",x"63",x"6F",x"6E", -- 0x3C38
    x"74",x"72",x"69",x"62",x"75",x"74",x"6F",x"72", -- 0x3C40
    x"73",x"20",x"74",x"6F",x"20",x"74",x"68",x"65", -- 0x3C48
    x"20",x"64",x"65",x"76",x"65",x"6C",x"6F",x"70", -- 0x3C50
    x"6D",x"65",x"6E",x"74",x"20",x"6F",x"66",x"20", -- 0x3C58
    x"74",x"68",x"65",x"20",x"42",x"42",x"43",x"20", -- 0x3C60
    x"43",x"6F",x"6D",x"70",x"75",x"74",x"65",x"72", -- 0x3C68
    x"20",x"28",x"61",x"6D",x"6F",x"6E",x"67",x"20", -- 0x3C70
    x"6F",x"74",x"68",x"65",x"72",x"73",x"20",x"74", -- 0x3C78
    x"6F",x"6F",x"20",x"6E",x"75",x"6D",x"65",x"72", -- 0x3C80
    x"6F",x"75",x"73",x"20",x"74",x"6F",x"20",x"6D", -- 0x3C88
    x"65",x"6E",x"74",x"69",x"6F",x"6E",x"29",x"3A", -- 0x3C90
    x"2D",x"20",x"44",x"61",x"76",x"69",x"64",x"20", -- 0x3C98
    x"41",x"6C",x"6C",x"65",x"6E",x"2C",x"42",x"6F", -- 0x3CA0
    x"62",x"20",x"41",x"75",x"73",x"74",x"69",x"6E", -- 0x3CA8
    x"2C",x"52",x"61",x"6D",x"20",x"42",x"61",x"6E", -- 0x3CB0
    x"65",x"72",x"6A",x"65",x"65",x"2C",x"50",x"61", -- 0x3CB8
    x"75",x"6C",x"20",x"42",x"6F",x"6E",x"64",x"2C", -- 0x3CC0
    x"41",x"6C",x"6C",x"65",x"6E",x"20",x"42",x"6F", -- 0x3CC8
    x"6F",x"74",x"68",x"72",x"6F",x"79",x"64",x"2C", -- 0x3CD0
    x"43",x"61",x"6D",x"62",x"72",x"69",x"64",x"67", -- 0x3CD8
    x"65",x"2C",x"43",x"6C",x"65",x"61",x"72",x"74", -- 0x3CE0
    x"6F",x"6E",x"65",x"2C",x"4A",x"6F",x"68",x"6E", -- 0x3CE8
    x"20",x"43",x"6F",x"6C",x"6C",x"2C",x"4A",x"6F", -- 0x3CF0
    x"68",x"6E",x"20",x"43",x"6F",x"78",x"2C",x"41", -- 0x3CF8
    x"6E",x"64",x"79",x"20",x"43",x"72",x"69",x"70", -- 0x3D00
    x"70",x"73",x"2C",x"43",x"68",x"72",x"69",x"73", -- 0x3D08
    x"20",x"43",x"75",x"72",x"72",x"79",x"2C",x"36", -- 0x3D10
    x"35",x"30",x"32",x"20",x"64",x"65",x"73",x"69", -- 0x3D18
    x"67",x"6E",x"65",x"72",x"73",x"2C",x"4A",x"65", -- 0x3D20
    x"72",x"65",x"6D",x"79",x"20",x"44",x"69",x"6F", -- 0x3D28
    x"6E",x"2C",x"54",x"69",x"6D",x"20",x"44",x"6F", -- 0x3D30
    x"62",x"73",x"6F",x"6E",x"2C",x"4A",x"6F",x"65", -- 0x3D38
    x"20",x"44",x"75",x"6E",x"6E",x"2C",x"50",x"61", -- 0x3D40
    x"75",x"6C",x"20",x"46",x"61",x"72",x"72",x"65", -- 0x3D48
    x"6C",x"6C",x"2C",x"46",x"65",x"72",x"72",x"61", -- 0x3D50
    x"6E",x"74",x"69",x"2C",x"53",x"74",x"65",x"76", -- 0x3D58
    x"65",x"20",x"46",x"75",x"72",x"62",x"65",x"72", -- 0x3D60
    x"2C",x"4A",x"6F",x"6E",x"20",x"47",x"69",x"62", -- 0x3D68
    x"62",x"6F",x"6E",x"73",x"2C",x"41",x"6E",x"64", -- 0x3D70
    x"72",x"65",x"77",x"20",x"47",x"6F",x"72",x"64", -- 0x3D78
    x"6F",x"6E",x"2C",x"4C",x"61",x"77",x"72",x"65", -- 0x3D80
    x"6E",x"63",x"65",x"20",x"48",x"61",x"72",x"64", -- 0x3D88
    x"77",x"69",x"63",x"6B",x"2C",x"44",x"79",x"6C", -- 0x3D90
    x"61",x"6E",x"20",x"48",x"61",x"72",x"72",x"69", -- 0x3D98
    x"73",x"2C",x"48",x"65",x"72",x"6D",x"61",x"6E", -- 0x3DA0
    x"6E",x"20",x"48",x"61",x"75",x"73",x"65",x"72", -- 0x3DA8
    x"2C",x"48",x"69",x"74",x"61",x"63",x"68",x"69", -- 0x3DB0
    x"2C",x"41",x"6E",x"64",x"79",x"20",x"48",x"6F", -- 0x3DB8
    x"70",x"70",x"65",x"72",x"2C",x"49",x"43",x"4C", -- 0x3DC0
    x"2C",x"4D",x"61",x"72",x"74",x"69",x"6E",x"20", -- 0x3DC8
    x"4A",x"61",x"63",x"6B",x"73",x"6F",x"6E",x"2C", -- 0x3DD0
    x"42",x"72",x"69",x"61",x"6E",x"20",x"4A",x"6F", -- 0x3DD8
    x"6E",x"65",x"73",x"2C",x"43",x"68",x"72",x"69", -- 0x3DE0
    x"73",x"20",x"4A",x"6F",x"72",x"64",x"61",x"6E", -- 0x3DE8
    x"2C",x"44",x"61",x"76",x"69",x"64",x"20",x"4B", -- 0x3DF0
    x"69",x"6E",x"67",x"2C",x"44",x"61",x"76",x"69", -- 0x3DF8
    x"64",x"20",x"4B",x"69",x"74",x"73",x"6F",x"6E", -- 0x3E00
    x"2C",x"50",x"61",x"75",x"6C",x"20",x"4B",x"72", -- 0x3E08
    x"69",x"77",x"61",x"63",x"7A",x"65",x"6B",x"2C", -- 0x3E10
    x"43",x"6F",x"6D",x"70",x"75",x"74",x"65",x"72", -- 0x3E18
    x"20",x"4C",x"61",x"62",x"6F",x"72",x"61",x"74", -- 0x3E20
    x"6F",x"72",x"79",x"2C",x"50",x"65",x"74",x"65", -- 0x3E28
    x"72",x"20",x"4D",x"69",x"6C",x"6C",x"65",x"72", -- 0x3E30
    x"2C",x"41",x"72",x"74",x"68",x"75",x"72",x"20", -- 0x3E38
    x"4E",x"6F",x"72",x"6D",x"61",x"6E",x"2C",x"47", -- 0x3E40
    x"6C",x"79",x"6E",x"20",x"50",x"68",x"69",x"6C", -- 0x3E48
    x"6C",x"69",x"70",x"73",x"2C",x"4D",x"69",x"6B", -- 0x3E50
    x"65",x"20",x"50",x"72",x"65",x"65",x"73",x"2C", -- 0x3E58
    x"4A",x"6F",x"68",x"6E",x"20",x"52",x"61",x"64", -- 0x3E60
    x"63",x"6C",x"69",x"66",x"66",x"65",x"2C",x"57", -- 0x3E68
    x"69",x"6C",x"62",x"65",x"72",x"66",x"6F",x"72", -- 0x3E70
    x"63",x"65",x"20",x"52",x"6F",x"61",x"64",x"2C", -- 0x3E78
    x"50",x"65",x"74",x"65",x"72",x"20",x"52",x"6F", -- 0x3E80
    x"62",x"69",x"6E",x"73",x"6F",x"6E",x"2C",x"52", -- 0x3E88
    x"69",x"63",x"68",x"61",x"72",x"64",x"20",x"52", -- 0x3E90
    x"75",x"73",x"73",x"65",x"6C",x"6C",x"2C",x"4B", -- 0x3E98
    x"69",x"6D",x"20",x"53",x"70",x"65",x"6E",x"63", -- 0x3EA0
    x"65",x"2D",x"4A",x"6F",x"6E",x"65",x"73",x"2C", -- 0x3EA8
    x"47",x"72",x"61",x"68",x"61",x"6D",x"20",x"54", -- 0x3EB0
    x"65",x"62",x"62",x"79",x"2C",x"4A",x"6F",x"6E", -- 0x3EB8
    x"20",x"54",x"68",x"61",x"63",x"6B",x"72",x"61", -- 0x3EC0
    x"79",x"2C",x"43",x"68",x"72",x"69",x"73",x"20", -- 0x3EC8
    x"54",x"75",x"72",x"6E",x"65",x"72",x"2C",x"41", -- 0x3ED0
    x"64",x"72",x"69",x"61",x"6E",x"20",x"57",x"61", -- 0x3ED8
    x"72",x"6E",x"65",x"72",x"2C",x"52",x"6F",x"67", -- 0x3EE0
    x"65",x"72",x"20",x"57",x"69",x"6C",x"73",x"6F", -- 0x3EE8
    x"6E",x"2C",x"41",x"6C",x"61",x"6E",x"20",x"57", -- 0x3EF0
    x"72",x"69",x"67",x"68",x"74",x"2E",x"CD",x"D9", -- 0x3EF8
    x"20",x"51",x"FF",x"20",x"51",x"FF",x"20",x"51", -- 0x3F00
    x"FF",x"20",x"51",x"FF",x"20",x"51",x"FF",x"20", -- 0x3F08
    x"51",x"FF",x"20",x"51",x"FF",x"20",x"51",x"FF", -- 0x3F10
    x"20",x"51",x"FF",x"20",x"51",x"FF",x"20",x"51", -- 0x3F18
    x"FF",x"20",x"51",x"FF",x"20",x"51",x"FF",x"20", -- 0x3F20
    x"51",x"FF",x"20",x"51",x"FF",x"20",x"51",x"FF", -- 0x3F28
    x"20",x"51",x"FF",x"20",x"51",x"FF",x"20",x"51", -- 0x3F30
    x"FF",x"20",x"51",x"FF",x"20",x"51",x"FF",x"20", -- 0x3F38
    x"51",x"FF",x"20",x"51",x"FF",x"20",x"51",x"FF", -- 0x3F40
    x"20",x"51",x"FF",x"20",x"51",x"FF",x"20",x"51", -- 0x3F48
    x"FF",x"48",x"48",x"48",x"48",x"48",x"08",x"48", -- 0x3F50
    x"8A",x"48",x"98",x"48",x"BA",x"A9",x"FF",x"9D", -- 0x3F58
    x"08",x"01",x"A9",x"88",x"9D",x"07",x"01",x"BC", -- 0x3F60
    x"0A",x"01",x"B9",x"9D",x"0D",x"9D",x"05",x"01", -- 0x3F68
    x"B9",x"9E",x"0D",x"9D",x"06",x"01",x"A5",x"F4", -- 0x3F70
    x"9D",x"09",x"01",x"B9",x"9F",x"0D",x"85",x"F4", -- 0x3F78
    x"8D",x"30",x"FE",x"68",x"A8",x"68",x"AA",x"68", -- 0x3F80
    x"40",x"08",x"48",x"8A",x"48",x"BA",x"BD",x"02", -- 0x3F88
    x"01",x"9D",x"05",x"01",x"BD",x"03",x"01",x"9D", -- 0x3F90
    x"06",x"01",x"68",x"AA",x"68",x"68",x"68",x"85", -- 0x3F98
    x"F4",x"8D",x"30",x"FE",x"68",x"28",x"60",x"8A", -- 0x3FA0
    x"B0",x"2A",x"BC",x"00",x"FC",x"60",x"BC",x"00", -- 0x3FA8
    x"FD",x"60",x"BC",x"00",x"FE",x"60",x"36",x"40", -- 0x3FB0
    x"D9",x"4C",x"0B",x"DC",x"4C",x"C0",x"C4",x"4C", -- 0x3FB8
    x"94",x"E4",x"4C",x"1E",x"EA",x"4C",x"2F",x"EA", -- 0x3FC0
    x"4C",x"C5",x"DE",x"4C",x"A4",x"E0",x"6C",x"1C", -- 0x3FC8
    x"02",x"6C",x"1A",x"02",x"6C",x"18",x"02",x"6C", -- 0x3FD0
    x"16",x"02",x"6C",x"14",x"02",x"6C",x"12",x"02", -- 0x3FD8
    x"6C",x"10",x"02",x"C9",x"0D",x"D0",x"07",x"A9", -- 0x3FE0
    x"0A",x"20",x"EE",x"FF",x"A9",x"0D",x"6C",x"0E", -- 0x3FE8
    x"02",x"6C",x"0C",x"02",x"6C",x"0A",x"02",x"6C", -- 0x3FF0
    x"08",x"02",x"00",x"0D",x"CD",x"D9",x"1C",x"DC"  -- 0x3FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
     DATA <= ROM(to_integer(unsigned(ADDR)));
  end process;
end RTL;
