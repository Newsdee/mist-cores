-- Copyright (C) 1991-2014 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.1.4 Build 182 03/12/2014 SJ Web Edition"
-- CREATED		"Thu Jul 10 07:36:50 2014"


LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY RS232 IS 
	PORT
	(
		store :  IN  STD_LOGIC;
		CTS :  IN  STD_LOGIC;
		Baudx4 :  IN  STD_LOGIC;
		RxD :  IN  STD_LOGIC;
		read :  IN  STD_LOGIC;
		i :  IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		TxD :  OUT  STD_LOGIC;
		RDY :  OUT  STD_LOGIC;
		snext :  OUT  STD_LOGIC;
		RTS :  OUT  STD_LOGIC;
		Y :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END RS232;

ARCHITECTURE bdf_type OF RS232 IS 

SIGNAL	Y_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	DFF_11 :  STD_LOGIC;
SIGNAL	DFF_124 :  STD_LOGIC;
SIGNAL	TFF_238 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	DFF_263 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	TFF_237 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	DFFE_inst :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;


BEGIN 
RDY <= DFF_11;
RTS <= DFF_263;
SYNTHESIZED_WIRE_22 <= '0';
SYNTHESIZED_WIRE_31 <= '1';
SYNTHESIZED_WIRE_34 <= '0';



PROCESS(SYNTHESIZED_WIRE_46,read)
BEGIN
IF (read = '0') THEN
	SYNTHESIZED_WIRE_48 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_46)) THEN
	SYNTHESIZED_WIRE_48 <= SYNTHESIZED_WIRE_47;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_46,read)
BEGIN
IF (read = '0') THEN
	DFF_11 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_46)) THEN
	DFF_11 <= SYNTHESIZED_WIRE_48;
END IF;
END PROCESS;


PROCESS(Baudx4,read)
BEGIN
IF (read = '0') THEN
	SYNTHESIZED_WIRE_49 <= '1';
ELSIF (RISING_EDGE(Baudx4)) THEN
	SYNTHESIZED_WIRE_49 <= SYNTHESIZED_WIRE_0;
END IF;
END PROCESS;


PROCESS(Baudx4,read)
BEGIN
IF (read = '0') THEN
	SYNTHESIZED_WIRE_46 <= '1';
ELSIF (RISING_EDGE(Baudx4)) THEN
	SYNTHESIZED_WIRE_46 <= SYNTHESIZED_WIRE_49;
END IF;
END PROCESS;


PROCESS(Baudx4,read)
BEGIN
IF (read = '0') THEN
	DFF_124 <= '1';
ELSIF (RISING_EDGE(Baudx4)) THEN
	DFF_124 <= SYNTHESIZED_WIRE_46;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_0 <= NOT(SYNTHESIZED_WIRE_50 AND DFF_11 AND DFF_124 AND SYNTHESIZED_WIRE_50 AND SYNTHESIZED_WIRE_46 AND SYNTHESIZED_WIRE_49);


SYNTHESIZED_WIRE_8 <= NOT(RxD);



PROCESS(Baudx4,SYNTHESIZED_WIRE_51)
BEGIN
IF (SYNTHESIZED_WIRE_51 = '0') THEN
	SYNTHESIZED_WIRE_52 <= '1';
ELSIF (RISING_EDGE(Baudx4)) THEN
	SYNTHESIZED_WIRE_52 <= TFF_238;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_52,SYNTHESIZED_WIRE_4,SYNTHESIZED_WIRE_5)
BEGIN
IF (SYNTHESIZED_WIRE_4 = '0') THEN
	SYNTHESIZED_WIRE_54 <= '0';
ELSIF (SYNTHESIZED_WIRE_5 = '0') THEN
	SYNTHESIZED_WIRE_54 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_52)) THEN
	SYNTHESIZED_WIRE_54 <= SYNTHESIZED_WIRE_53;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_52,SYNTHESIZED_WIRE_6,SYNTHESIZED_WIRE_7)
BEGIN
IF (SYNTHESIZED_WIRE_6 = '0') THEN
	SYNTHESIZED_WIRE_55 <= '0';
ELSIF (SYNTHESIZED_WIRE_7 = '0') THEN
	SYNTHESIZED_WIRE_55 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_52)) THEN
	SYNTHESIZED_WIRE_55 <= SYNTHESIZED_WIRE_54;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_52,store)
BEGIN
IF (store = '0') THEN
	SYNTHESIZED_WIRE_56 <= '0';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_52)) THEN
	SYNTHESIZED_WIRE_56 <= SYNTHESIZED_WIRE_55;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_50 <= SYNTHESIZED_WIRE_8 OR DFF_263;


PROCESS(SYNTHESIZED_WIRE_52,SYNTHESIZED_WIRE_9)
BEGIN
IF (SYNTHESIZED_WIRE_9 = '0') THEN
	TxD <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_52)) THEN
	TxD <= SYNTHESIZED_WIRE_56;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_52,SYNTHESIZED_WIRE_10,SYNTHESIZED_WIRE_11)
BEGIN
IF (SYNTHESIZED_WIRE_10 = '0') THEN
	SYNTHESIZED_WIRE_53 <= '0';
ELSIF (SYNTHESIZED_WIRE_11 = '0') THEN
	SYNTHESIZED_WIRE_53 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_52)) THEN
	SYNTHESIZED_WIRE_53 <= SYNTHESIZED_WIRE_57;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_52,SYNTHESIZED_WIRE_12,SYNTHESIZED_WIRE_13)
BEGIN
IF (SYNTHESIZED_WIRE_12 = '0') THEN
	SYNTHESIZED_WIRE_57 <= '0';
ELSIF (SYNTHESIZED_WIRE_13 = '0') THEN
	SYNTHESIZED_WIRE_57 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_52)) THEN
	SYNTHESIZED_WIRE_57 <= SYNTHESIZED_WIRE_58;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_52,SYNTHESIZED_WIRE_14,SYNTHESIZED_WIRE_15)
BEGIN
IF (SYNTHESIZED_WIRE_14 = '0') THEN
	SYNTHESIZED_WIRE_58 <= '0';
ELSIF (SYNTHESIZED_WIRE_15 = '0') THEN
	SYNTHESIZED_WIRE_58 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_52)) THEN
	SYNTHESIZED_WIRE_58 <= SYNTHESIZED_WIRE_59;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_52,SYNTHESIZED_WIRE_16,SYNTHESIZED_WIRE_17)
BEGIN
IF (SYNTHESIZED_WIRE_16 = '0') THEN
	SYNTHESIZED_WIRE_59 <= '0';
ELSIF (SYNTHESIZED_WIRE_17 = '0') THEN
	SYNTHESIZED_WIRE_59 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_52)) THEN
	SYNTHESIZED_WIRE_59 <= SYNTHESIZED_WIRE_60;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_52,SYNTHESIZED_WIRE_18,SYNTHESIZED_WIRE_19)
BEGIN
IF (SYNTHESIZED_WIRE_18 = '0') THEN
	SYNTHESIZED_WIRE_60 <= '0';
ELSIF (SYNTHESIZED_WIRE_19 = '0') THEN
	SYNTHESIZED_WIRE_60 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_52)) THEN
	SYNTHESIZED_WIRE_60 <= SYNTHESIZED_WIRE_61;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_52,SYNTHESIZED_WIRE_20,SYNTHESIZED_WIRE_21)
BEGIN
IF (SYNTHESIZED_WIRE_20 = '0') THEN
	SYNTHESIZED_WIRE_61 <= '0';
ELSIF (SYNTHESIZED_WIRE_21 = '0') THEN
	SYNTHESIZED_WIRE_61 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_52)) THEN
	SYNTHESIZED_WIRE_61 <= SYNTHESIZED_WIRE_62;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_52,store)
BEGIN
IF (store = '0') THEN
	SYNTHESIZED_WIRE_62 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_52)) THEN
	SYNTHESIZED_WIRE_62 <= SYNTHESIZED_WIRE_22;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_19 <= NOT(SYNTHESIZED_WIRE_63 AND i(6));


SYNTHESIZED_WIRE_21 <= NOT(SYNTHESIZED_WIRE_63 AND i(7));


SYNTHESIZED_WIRE_18 <= i(6) OR store;


SYNTHESIZED_WIRE_20 <= i(7) OR store;


SYNTHESIZED_WIRE_15 <= NOT(SYNTHESIZED_WIRE_63 AND i(4));


SYNTHESIZED_WIRE_17 <= NOT(SYNTHESIZED_WIRE_63 AND i(5));


SYNTHESIZED_WIRE_14 <= i(4) OR store;


SYNTHESIZED_WIRE_16 <= i(5) OR store;


SYNTHESIZED_WIRE_11 <= NOT(SYNTHESIZED_WIRE_63 AND i(2));


SYNTHESIZED_WIRE_13 <= NOT(SYNTHESIZED_WIRE_63 AND i(3));


SYNTHESIZED_WIRE_10 <= i(2) OR store;


SYNTHESIZED_WIRE_12 <= i(3) OR store;


SYNTHESIZED_WIRE_5 <= NOT(SYNTHESIZED_WIRE_63 AND i(1));


SYNTHESIZED_WIRE_4 <= i(1) OR store;



SYNTHESIZED_WIRE_7 <= NOT(SYNTHESIZED_WIRE_63 AND i(0));


SYNTHESIZED_WIRE_6 <= i(0) OR store;


SYNTHESIZED_WIRE_32 <= SYNTHESIZED_WIRE_56 OR SYNTHESIZED_WIRE_55 OR SYNTHESIZED_WIRE_54 OR SYNTHESIZED_WIRE_53 OR SYNTHESIZED_WIRE_57 OR SYNTHESIZED_WIRE_58 OR SYNTHESIZED_WIRE_59 OR SYNTHESIZED_WIRE_60;


SYNTHESIZED_WIRE_63 <= NOT(store);



PROCESS(Baudx4)
VARIABLE TFF_237_synthesized_var : STD_LOGIC;
BEGIN
IF (RISING_EDGE(Baudx4)) THEN
	TFF_237_synthesized_var := TFF_237_synthesized_var XOR SYNTHESIZED_WIRE_31;
END IF;
	TFF_237 <= TFF_237_synthesized_var;
END PROCESS;


PROCESS(Baudx4)
VARIABLE TFF_238_synthesized_var : STD_LOGIC;
BEGIN
IF (RISING_EDGE(Baudx4)) THEN
	TFF_238_synthesized_var := TFF_238_synthesized_var XOR TFF_237;
END IF;
	TFF_238 <= TFF_238_synthesized_var;
END PROCESS;



SYNTHESIZED_WIRE_51 <= SYNTHESIZED_WIRE_32 OR SYNTHESIZED_WIRE_62 OR SYNTHESIZED_WIRE_61;


SYNTHESIZED_WIRE_9 <= store AND SYNTHESIZED_WIRE_51;


PROCESS(read,SYNTHESIZED_WIRE_46)
BEGIN
IF (SYNTHESIZED_WIRE_46 = '0') THEN
	DFF_263 <= '1';
ELSIF (RISING_EDGE(read)) THEN
	DFF_263 <= SYNTHESIZED_WIRE_34;
END IF;
END PROCESS;



SYNTHESIZED_WIRE_45 <= NOT(SYNTHESIZED_WIRE_48);



PROCESS(SYNTHESIZED_WIRE_46,read)
BEGIN
IF (read = '0') THEN
	SYNTHESIZED_WIRE_64 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_46)) THEN
	SYNTHESIZED_WIRE_64 <= RxD;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_46,read)
BEGIN
IF (read = '0') THEN
	SYNTHESIZED_WIRE_65 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_46)) THEN
	SYNTHESIZED_WIRE_65 <= SYNTHESIZED_WIRE_64;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_46,read)
BEGIN
IF (read = '0') THEN
	SYNTHESIZED_WIRE_66 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_46)) THEN
	SYNTHESIZED_WIRE_66 <= SYNTHESIZED_WIRE_65;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_46,read)
BEGIN
IF (read = '0') THEN
	SYNTHESIZED_WIRE_67 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_46)) THEN
	SYNTHESIZED_WIRE_67 <= SYNTHESIZED_WIRE_66;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_46,read)
BEGIN
IF (read = '0') THEN
	SYNTHESIZED_WIRE_68 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_46)) THEN
	SYNTHESIZED_WIRE_68 <= SYNTHESIZED_WIRE_67;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_46,read)
BEGIN
IF (read = '0') THEN
	SYNTHESIZED_WIRE_69 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_46)) THEN
	SYNTHESIZED_WIRE_69 <= SYNTHESIZED_WIRE_68;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_46,read)
BEGIN
IF (read = '0') THEN
	SYNTHESIZED_WIRE_47 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_46)) THEN
	SYNTHESIZED_WIRE_47 <= SYNTHESIZED_WIRE_69;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_46,read)
BEGIN
IF (read = '0') THEN
	DFFE_inst <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_46)) THEN
	IF (SYNTHESIZED_WIRE_70 = '1') THEN
	DFFE_inst <= SYNTHESIZED_WIRE_48;
	END IF;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_46)
BEGIN
IF (RISING_EDGE(SYNTHESIZED_WIRE_46)) THEN
	IF (SYNTHESIZED_WIRE_70 = '1') THEN
	Y_ALTERA_SYNTHESIZED(0) <= SYNTHESIZED_WIRE_47;
	END IF;
END IF;
END PROCESS;


snext <= NOT(SYNTHESIZED_WIRE_51 OR CTS);


PROCESS(SYNTHESIZED_WIRE_46)
BEGIN
IF (RISING_EDGE(SYNTHESIZED_WIRE_46)) THEN
	IF (SYNTHESIZED_WIRE_70 = '1') THEN
	Y_ALTERA_SYNTHESIZED(1) <= SYNTHESIZED_WIRE_69;
	END IF;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_46)
BEGIN
IF (RISING_EDGE(SYNTHESIZED_WIRE_46)) THEN
	IF (SYNTHESIZED_WIRE_70 = '1') THEN
	Y_ALTERA_SYNTHESIZED(2) <= SYNTHESIZED_WIRE_68;
	END IF;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_46)
BEGIN
IF (RISING_EDGE(SYNTHESIZED_WIRE_46)) THEN
	IF (SYNTHESIZED_WIRE_70 = '1') THEN
	Y_ALTERA_SYNTHESIZED(3) <= SYNTHESIZED_WIRE_67;
	END IF;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_46)
BEGIN
IF (RISING_EDGE(SYNTHESIZED_WIRE_46)) THEN
	IF (SYNTHESIZED_WIRE_70 = '1') THEN
	Y_ALTERA_SYNTHESIZED(4) <= SYNTHESIZED_WIRE_66;
	END IF;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_46)
BEGIN
IF (RISING_EDGE(SYNTHESIZED_WIRE_46)) THEN
	IF (SYNTHESIZED_WIRE_70 = '1') THEN
	Y_ALTERA_SYNTHESIZED(5) <= SYNTHESIZED_WIRE_65;
	END IF;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_46)
BEGIN
IF (RISING_EDGE(SYNTHESIZED_WIRE_46)) THEN
	IF (SYNTHESIZED_WIRE_70 = '1') THEN
	Y_ALTERA_SYNTHESIZED(6) <= SYNTHESIZED_WIRE_64;
	END IF;
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_46)
BEGIN
IF (RISING_EDGE(SYNTHESIZED_WIRE_46)) THEN
	IF (SYNTHESIZED_WIRE_70 = '1') THEN
	Y_ALTERA_SYNTHESIZED(7) <= RxD;
	END IF;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_70 <= DFFE_inst AND SYNTHESIZED_WIRE_45;

Y <= Y_ALTERA_SYNTHESIZED;

END bdf_type;